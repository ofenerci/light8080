//-----------------------------------------------------------------------------
//
// RAM image for input code file: hello.hex
//
//-----------------------------------------------------------------------------
module ram_image
(
	clk, addr, 
	we, din, dout
);
//-----------------------------------------------------------------------------
input           clk;
input   [11:0]  addr;
input           we;
input   [7:0]   din;
output  [7:0]   dout;
//-----------------------------------------------------------------------------
reg [7:0] dout;
reg [7:0] ram [4095:0];
//-----------------------------------------------------------------------------
initial 
begin
    ram[0] = 8'h21; ram[1] = 8'h00; ram[2] = 8'h0c; ram[3] = 8'hf9; 
    ram[4] = 8'hcd; ram[5] = 8'he3; ram[6] = 8'h02; ram[7] = 8'h7e; 
    ram[8] = 8'h6f; ram[9] = 8'h07; ram[10] = 8'h9f; ram[11] = 8'h67; 
    ram[12] = 8'hc9; ram[13] = 8'h7e; ram[14] = 8'h23; ram[15] = 8'h66; 
    ram[16] = 8'h6f; ram[17] = 8'hc9; ram[18] = 8'h7d; ram[19] = 8'h12; 
    ram[20] = 8'hc9; ram[21] = 8'h7d; ram[22] = 8'h12; ram[23] = 8'h13; 
    ram[24] = 8'h7c; ram[25] = 8'h12; ram[26] = 8'hc9; ram[27] = 8'h7d; 
    ram[28] = 8'hb3; ram[29] = 8'h6f; ram[30] = 8'h7c; ram[31] = 8'hb2; 
    ram[32] = 8'h67; ram[33] = 8'hc9; ram[34] = 8'h7d; ram[35] = 8'hab; 
    ram[36] = 8'h6f; ram[37] = 8'h7c; ram[38] = 8'haa; ram[39] = 8'h67; 
    ram[40] = 8'hc9; ram[41] = 8'h7d; ram[42] = 8'ha3; ram[43] = 8'h6f; 
    ram[44] = 8'h7c; ram[45] = 8'ha2; ram[46] = 8'h67; ram[47] = 8'hc9; 
    ram[48] = 8'hcd; ram[49] = 8'h56; ram[50] = 8'h00; ram[51] = 8'hc8; 
    ram[52] = 8'h2b; ram[53] = 8'hc9; ram[54] = 8'hcd; ram[55] = 8'h56; 
    ram[56] = 8'h00; ram[57] = 8'hc0; ram[58] = 8'h2b; ram[59] = 8'hc9; 
    ram[60] = 8'heb; ram[61] = 8'hcd; ram[62] = 8'h56; ram[63] = 8'h00; 
    ram[64] = 8'hd8; ram[65] = 8'h2b; ram[66] = 8'hc9; ram[67] = 8'hcd; 
    ram[68] = 8'h56; ram[69] = 8'h00; ram[70] = 8'hc8; ram[71] = 8'hd8; 
    ram[72] = 8'h2b; ram[73] = 8'hc9; ram[74] = 8'hcd; ram[75] = 8'h56; 
    ram[76] = 8'h00; ram[77] = 8'hd0; ram[78] = 8'h2b; ram[79] = 8'hc9; 
    ram[80] = 8'hcd; ram[81] = 8'h56; ram[82] = 8'h00; ram[83] = 8'hd8; 
    ram[84] = 8'h2b; ram[85] = 8'hc9; ram[86] = 8'h7b; ram[87] = 8'h95; 
    ram[88] = 8'h5f; ram[89] = 8'h7a; ram[90] = 8'h9c; ram[91] = 8'h21; 
    ram[92] = 8'h01; ram[93] = 8'h00; ram[94] = 8'hfa; ram[95] = 8'h63; 
    ram[96] = 8'h00; ram[97] = 8'hb3; ram[98] = 8'hc9; ram[99] = 8'hb3; 
    ram[100] = 8'h37; ram[101] = 8'hc9; ram[102] = 8'hcd; ram[103] = 8'h80; 
    ram[104] = 8'h00; ram[105] = 8'hd0; ram[106] = 8'h2b; ram[107] = 8'hc9; 
    ram[108] = 8'hcd; ram[109] = 8'h80; ram[110] = 8'h00; ram[111] = 8'hd8; 
    ram[112] = 8'h2b; ram[113] = 8'hc9; ram[114] = 8'heb; ram[115] = 8'hcd; 
    ram[116] = 8'h80; ram[117] = 8'h00; ram[118] = 8'hd8; ram[119] = 8'h2b; 
    ram[120] = 8'hc9; ram[121] = 8'hcd; ram[122] = 8'h80; ram[123] = 8'h00; 
    ram[124] = 8'hc8; ram[125] = 8'hd8; ram[126] = 8'h2b; ram[127] = 8'hc9; 
    ram[128] = 8'h7a; ram[129] = 8'hbc; ram[130] = 8'hc2; ram[131] = 8'h87; 
    ram[132] = 8'h00; ram[133] = 8'h7b; ram[134] = 8'hbd; ram[135] = 8'h21; 
    ram[136] = 8'h01; ram[137] = 8'h00; ram[138] = 8'hc9; ram[139] = 8'heb; 
    ram[140] = 8'h7c; ram[141] = 8'h17; ram[142] = 8'h7c; ram[143] = 8'h1f; 
    ram[144] = 8'h67; ram[145] = 8'h7d; ram[146] = 8'h1f; ram[147] = 8'h6f; 
    ram[148] = 8'h1d; ram[149] = 8'hc2; ram[150] = 8'h8c; ram[151] = 8'h00; 
    ram[152] = 8'hc9; ram[153] = 8'heb; ram[154] = 8'h29; ram[155] = 8'h1d; 
    ram[156] = 8'hc2; ram[157] = 8'h9a; ram[158] = 8'h00; ram[159] = 8'hc9; 
    ram[160] = 8'h7b; ram[161] = 8'h95; ram[162] = 8'h6f; ram[163] = 8'h7a; 
    ram[164] = 8'h9c; ram[165] = 8'h67; ram[166] = 8'hc9; ram[167] = 8'hcd; 
    ram[168] = 8'hac; ram[169] = 8'h00; ram[170] = 8'h23; ram[171] = 8'hc9; 
    ram[172] = 8'h7c; ram[173] = 8'h2f; ram[174] = 8'h67; ram[175] = 8'h7d; 
    ram[176] = 8'h2f; ram[177] = 8'h6f; ram[178] = 8'hc9; ram[179] = 8'h44; 
    ram[180] = 8'h4d; ram[181] = 8'h21; ram[182] = 8'h00; ram[183] = 8'h00; 
    ram[184] = 8'h79; ram[185] = 8'h0f; ram[186] = 8'hd2; ram[187] = 8'hbe; 
    ram[188] = 8'h00; ram[189] = 8'h19; ram[190] = 8'haf; ram[191] = 8'h78; 
    ram[192] = 8'h1f; ram[193] = 8'h47; ram[194] = 8'h79; ram[195] = 8'h1f; 
    ram[196] = 8'h4f; ram[197] = 8'hb0; ram[198] = 8'hc8; ram[199] = 8'haf; 
    ram[200] = 8'h7b; ram[201] = 8'h17; ram[202] = 8'h5f; ram[203] = 8'h7a; 
    ram[204] = 8'h17; ram[205] = 8'h57; ram[206] = 8'hb3; ram[207] = 8'hc8; 
    ram[208] = 8'hc3; ram[209] = 8'hb8; ram[210] = 8'h00; ram[211] = 8'h44; 
    ram[212] = 8'h4d; ram[213] = 8'h7a; ram[214] = 8'ha8; ram[215] = 8'hf5; 
    ram[216] = 8'h7a; ram[217] = 8'hb7; ram[218] = 8'hfc; ram[219] = 8'h14; 
    ram[220] = 8'h01; ram[221] = 8'h78; ram[222] = 8'hb7; ram[223] = 8'hfc; 
    ram[224] = 8'h1c; ram[225] = 8'h01; ram[226] = 8'h3e; ram[227] = 8'h10; 
    ram[228] = 8'hf5; ram[229] = 8'heb; ram[230] = 8'h11; ram[231] = 8'h00; 
    ram[232] = 8'h00; ram[233] = 8'h29; ram[234] = 8'hcd; ram[235] = 8'h24; 
    ram[236] = 8'h01; ram[237] = 8'hca; ram[238] = 8'h00; ram[239] = 8'h01; 
    ram[240] = 8'hcd; ram[241] = 8'h2c; ram[242] = 8'h01; ram[243] = 8'hfa; 
    ram[244] = 8'h00; ram[245] = 8'h01; ram[246] = 8'h7d; ram[247] = 8'hf6; 
    ram[248] = 8'h01; ram[249] = 8'h6f; ram[250] = 8'h7b; ram[251] = 8'h91; 
    ram[252] = 8'h5f; ram[253] = 8'h7a; ram[254] = 8'h98; ram[255] = 8'h57; 
    ram[256] = 8'hf1; ram[257] = 8'h3d; ram[258] = 8'hca; ram[259] = 8'h09; 
    ram[260] = 8'h01; ram[261] = 8'hf5; ram[262] = 8'hc3; ram[263] = 8'he9; 
    ram[264] = 8'h00; ram[265] = 8'hf1; ram[266] = 8'hf0; ram[267] = 8'hcd; 
    ram[268] = 8'h14; ram[269] = 8'h01; ram[270] = 8'heb; ram[271] = 8'hcd; 
    ram[272] = 8'h14; ram[273] = 8'h01; ram[274] = 8'heb; ram[275] = 8'hc9; 
    ram[276] = 8'h7a; ram[277] = 8'h2f; ram[278] = 8'h57; ram[279] = 8'h7b; 
    ram[280] = 8'h2f; ram[281] = 8'h5f; ram[282] = 8'h13; ram[283] = 8'hc9; 
    ram[284] = 8'h78; ram[285] = 8'h2f; ram[286] = 8'h47; ram[287] = 8'h79; 
    ram[288] = 8'h2f; ram[289] = 8'h4f; ram[290] = 8'h03; ram[291] = 8'hc9; 
    ram[292] = 8'h7b; ram[293] = 8'h17; ram[294] = 8'h5f; ram[295] = 8'h7a; 
    ram[296] = 8'h17; ram[297] = 8'h57; ram[298] = 8'hb3; ram[299] = 8'hc9; 
    ram[300] = 8'h7b; ram[301] = 8'h91; ram[302] = 8'h7a; ram[303] = 8'h98; 
    ram[304] = 8'hc9; ram[305] = 8'hdb; ram[306] = 8'h83; ram[307] = 8'hcf; 
    ram[308] = 8'he5; ram[309] = 8'h21; ram[310] = 8'h01; ram[311] = 8'h00; 
    ram[312] = 8'hd1; ram[313] = 8'hcd; ram[314] = 8'h29; ram[315] = 8'h00; 
    ram[316] = 8'h7c; ram[317] = 8'hb5; ram[318] = 8'hca; ram[319] = 8'h44; 
    ram[320] = 8'h01; ram[321] = 8'hc3; ram[322] = 8'h31; ram[323] = 8'h01; 
    ram[324] = 8'h21; ram[325] = 8'h02; ram[326] = 8'h00; ram[327] = 8'h39; 
    ram[328] = 8'hcd; ram[329] = 8'h07; ram[330] = 8'h00; ram[331] = 8'h7d; 
    ram[332] = 8'hd3; ram[333] = 8'h80; ram[334] = 8'hc9; ram[335] = 8'hdb; 
    ram[336] = 8'h83; ram[337] = 8'hcf; ram[338] = 8'he5; ram[339] = 8'h21; 
    ram[340] = 8'h10; ram[341] = 8'h00; ram[342] = 8'hd1; ram[343] = 8'hcd; 
    ram[344] = 8'h29; ram[345] = 8'h00; ram[346] = 8'h7c; ram[347] = 8'hb5; 
    ram[348] = 8'hca; ram[349] = 8'h6d; ram[350] = 8'h01; ram[351] = 8'hdb; 
    ram[352] = 8'h80; ram[353] = 8'hcf; ram[354] = 8'h7d; ram[355] = 8'h32; 
    ram[356] = 8'h9e; ram[357] = 8'h03; ram[358] = 8'h21; ram[359] = 8'h01; 
    ram[360] = 8'h00; ram[361] = 8'hc9; ram[362] = 8'hc3; ram[363] = 8'h71; 
    ram[364] = 8'h01; ram[365] = 8'h21; ram[366] = 8'h00; ram[367] = 8'h00; 
    ram[368] = 8'hc9; ram[369] = 8'hc9; ram[370] = 8'h21; ram[371] = 8'h0d; 
    ram[372] = 8'h00; ram[373] = 8'he5; ram[374] = 8'hcd; ram[375] = 8'h31; 
    ram[376] = 8'h01; ram[377] = 8'hc1; ram[378] = 8'h21; ram[379] = 8'h0a; 
    ram[380] = 8'h00; ram[381] = 8'he5; ram[382] = 8'hcd; ram[383] = 8'h31; 
    ram[384] = 8'h01; ram[385] = 8'hc1; ram[386] = 8'hc9; ram[387] = 8'h21; 
    ram[388] = 8'h02; ram[389] = 8'h00; ram[390] = 8'h39; ram[391] = 8'hcd; 
    ram[392] = 8'h0d; ram[393] = 8'h00; ram[394] = 8'hcd; ram[395] = 8'h07; 
    ram[396] = 8'h00; ram[397] = 8'he5; ram[398] = 8'h21; ram[399] = 8'h00; 
    ram[400] = 8'h00; ram[401] = 8'hd1; ram[402] = 8'hcd; ram[403] = 8'h36; 
    ram[404] = 8'h00; ram[405] = 8'h7c; ram[406] = 8'hb5; ram[407] = 8'hca; 
    ram[408] = 8'hb3; ram[409] = 8'h01; ram[410] = 8'h21; ram[411] = 8'h02; 
    ram[412] = 8'h00; ram[413] = 8'h39; ram[414] = 8'he5; ram[415] = 8'hcd; 
    ram[416] = 8'h0d; ram[417] = 8'h00; ram[418] = 8'h23; ram[419] = 8'hd1; 
    ram[420] = 8'hcd; ram[421] = 8'h15; ram[422] = 8'h00; ram[423] = 8'h2b; 
    ram[424] = 8'hcd; ram[425] = 8'h07; ram[426] = 8'h00; ram[427] = 8'he5; 
    ram[428] = 8'hcd; ram[429] = 8'h31; ram[430] = 8'h01; ram[431] = 8'hc1; 
    ram[432] = 8'hc3; ram[433] = 8'h83; ram[434] = 8'h01; ram[435] = 8'hc9; 
    ram[436] = 8'h21; ram[437] = 8'h02; ram[438] = 8'h00; ram[439] = 8'h39; 
    ram[440] = 8'hcd; ram[441] = 8'h0d; ram[442] = 8'h00; ram[443] = 8'he5; 
    ram[444] = 8'h21; ram[445] = 8'h00; ram[446] = 8'h00; ram[447] = 8'hd1; 
    ram[448] = 8'hcd; ram[449] = 8'h50; ram[450] = 8'h00; ram[451] = 8'h7c; 
    ram[452] = 8'hb5; ram[453] = 8'hca; ram[454] = 8'he3; ram[455] = 8'h01; 
    ram[456] = 8'h21; ram[457] = 8'h2d; ram[458] = 8'h00; ram[459] = 8'he5; 
    ram[460] = 8'hcd; ram[461] = 8'h31; ram[462] = 8'h01; ram[463] = 8'hc1; 
    ram[464] = 8'h21; ram[465] = 8'h02; ram[466] = 8'h00; ram[467] = 8'h39; 
    ram[468] = 8'he5; ram[469] = 8'h21; ram[470] = 8'h04; ram[471] = 8'h00; 
    ram[472] = 8'h39; ram[473] = 8'hcd; ram[474] = 8'h0d; ram[475] = 8'h00; 
    ram[476] = 8'hcd; ram[477] = 8'ha7; ram[478] = 8'h00; ram[479] = 8'hd1; 
    ram[480] = 8'hcd; ram[481] = 8'h15; ram[482] = 8'h00; ram[483] = 8'h21; 
    ram[484] = 8'h02; ram[485] = 8'h00; ram[486] = 8'h39; ram[487] = 8'hcd; 
    ram[488] = 8'h0d; ram[489] = 8'h00; ram[490] = 8'he5; ram[491] = 8'hcd; 
    ram[492] = 8'hf0; ram[493] = 8'h01; ram[494] = 8'hc1; ram[495] = 8'hc9; 
    ram[496] = 8'hc5; ram[497] = 8'h21; ram[498] = 8'h00; ram[499] = 8'h00; 
    ram[500] = 8'h39; ram[501] = 8'he5; ram[502] = 8'h21; ram[503] = 8'h06; 
    ram[504] = 8'h00; ram[505] = 8'h39; ram[506] = 8'hcd; ram[507] = 8'h0d; 
    ram[508] = 8'h00; ram[509] = 8'he5; ram[510] = 8'h21; ram[511] = 8'h0a; 
    ram[512] = 8'h00; ram[513] = 8'hd1; ram[514] = 8'hcd; ram[515] = 8'hd3; 
    ram[516] = 8'h00; ram[517] = 8'hd1; ram[518] = 8'hcd; ram[519] = 8'h15; 
    ram[520] = 8'h00; ram[521] = 8'h21; ram[522] = 8'h00; ram[523] = 8'h00; 
    ram[524] = 8'h39; ram[525] = 8'hcd; ram[526] = 8'h0d; ram[527] = 8'h00; 
    ram[528] = 8'h7c; ram[529] = 8'hb5; ram[530] = 8'hca; ram[531] = 8'h21; 
    ram[532] = 8'h02; ram[533] = 8'h21; ram[534] = 8'h00; ram[535] = 8'h00; 
    ram[536] = 8'h39; ram[537] = 8'hcd; ram[538] = 8'h0d; ram[539] = 8'h00; 
    ram[540] = 8'he5; ram[541] = 8'hcd; ram[542] = 8'hf0; ram[543] = 8'h01; 
    ram[544] = 8'hc1; ram[545] = 8'h21; ram[546] = 8'h30; ram[547] = 8'h00; 
    ram[548] = 8'he5; ram[549] = 8'h21; ram[550] = 8'h06; ram[551] = 8'h00; 
    ram[552] = 8'h39; ram[553] = 8'hcd; ram[554] = 8'h0d; ram[555] = 8'h00; 
    ram[556] = 8'he5; ram[557] = 8'h21; ram[558] = 8'h04; ram[559] = 8'h00; 
    ram[560] = 8'h39; ram[561] = 8'hcd; ram[562] = 8'h0d; ram[563] = 8'h00; 
    ram[564] = 8'he5; ram[565] = 8'h21; ram[566] = 8'h0a; ram[567] = 8'h00; 
    ram[568] = 8'hd1; ram[569] = 8'hcd; ram[570] = 8'hb3; ram[571] = 8'h00; 
    ram[572] = 8'hd1; ram[573] = 8'hcd; ram[574] = 8'ha0; ram[575] = 8'h00; 
    ram[576] = 8'hd1; ram[577] = 8'h19; ram[578] = 8'he5; ram[579] = 8'hcd; 
    ram[580] = 8'h31; ram[581] = 8'h01; ram[582] = 8'hc1; ram[583] = 8'hc1; 
    ram[584] = 8'hc9; ram[585] = 8'hc5; ram[586] = 8'h21; ram[587] = 8'h00; 
    ram[588] = 8'h00; ram[589] = 8'h39; ram[590] = 8'he5; ram[591] = 8'h21; 
    ram[592] = 8'h06; ram[593] = 8'h00; ram[594] = 8'h39; ram[595] = 8'hcd; 
    ram[596] = 8'h0d; ram[597] = 8'h00; ram[598] = 8'he5; ram[599] = 8'h21; 
    ram[600] = 8'h10; ram[601] = 8'h00; ram[602] = 8'hd1; ram[603] = 8'hcd; 
    ram[604] = 8'hd3; ram[605] = 8'h00; ram[606] = 8'hd1; ram[607] = 8'hcd; 
    ram[608] = 8'h15; ram[609] = 8'h00; ram[610] = 8'h21; ram[611] = 8'h00; 
    ram[612] = 8'h00; ram[613] = 8'h39; ram[614] = 8'hcd; ram[615] = 8'h0d; 
    ram[616] = 8'h00; ram[617] = 8'h7c; ram[618] = 8'hb5; ram[619] = 8'hca; 
    ram[620] = 8'h7a; ram[621] = 8'h02; ram[622] = 8'h21; ram[623] = 8'h00; 
    ram[624] = 8'h00; ram[625] = 8'h39; ram[626] = 8'hcd; ram[627] = 8'h0d; 
    ram[628] = 8'h00; ram[629] = 8'he5; ram[630] = 8'hcd; ram[631] = 8'h49; 
    ram[632] = 8'h02; ram[633] = 8'hc1; ram[634] = 8'h21; ram[635] = 8'h00; 
    ram[636] = 8'h00; ram[637] = 8'h39; ram[638] = 8'he5; ram[639] = 8'h21; 
    ram[640] = 8'h06; ram[641] = 8'h00; ram[642] = 8'h39; ram[643] = 8'hcd; 
    ram[644] = 8'h0d; ram[645] = 8'h00; ram[646] = 8'he5; ram[647] = 8'h21; 
    ram[648] = 8'h04; ram[649] = 8'h00; ram[650] = 8'h39; ram[651] = 8'hcd; 
    ram[652] = 8'h0d; ram[653] = 8'h00; ram[654] = 8'he5; ram[655] = 8'h21; 
    ram[656] = 8'h10; ram[657] = 8'h00; ram[658] = 8'hd1; ram[659] = 8'hcd; 
    ram[660] = 8'hb3; ram[661] = 8'h00; ram[662] = 8'hd1; ram[663] = 8'hcd; 
    ram[664] = 8'ha0; ram[665] = 8'h00; ram[666] = 8'hd1; ram[667] = 8'hcd; 
    ram[668] = 8'h15; ram[669] = 8'h00; ram[670] = 8'h21; ram[671] = 8'h00; 
    ram[672] = 8'h00; ram[673] = 8'h39; ram[674] = 8'hcd; ram[675] = 8'h0d; 
    ram[676] = 8'h00; ram[677] = 8'he5; ram[678] = 8'h21; ram[679] = 8'h09; 
    ram[680] = 8'h00; ram[681] = 8'hd1; ram[682] = 8'hcd; ram[683] = 8'h3c; 
    ram[684] = 8'h00; ram[685] = 8'h7c; ram[686] = 8'hb5; ram[687] = 8'hca; 
    ram[688] = 8'hcf; ram[689] = 8'h02; ram[690] = 8'h21; ram[691] = 8'h41; 
    ram[692] = 8'h00; ram[693] = 8'he5; ram[694] = 8'h21; ram[695] = 8'h02; 
    ram[696] = 8'h00; ram[697] = 8'h39; ram[698] = 8'hcd; ram[699] = 8'h0d; 
    ram[700] = 8'h00; ram[701] = 8'hd1; ram[702] = 8'h19; ram[703] = 8'he5; 
    ram[704] = 8'h21; ram[705] = 8'h0a; ram[706] = 8'h00; ram[707] = 8'hd1; 
    ram[708] = 8'hcd; ram[709] = 8'ha0; ram[710] = 8'h00; ram[711] = 8'he5; 
    ram[712] = 8'hcd; ram[713] = 8'h31; ram[714] = 8'h01; ram[715] = 8'hc1; 
    ram[716] = 8'hc3; ram[717] = 8'he1; ram[718] = 8'h02; ram[719] = 8'h21; 
    ram[720] = 8'h30; ram[721] = 8'h00; ram[722] = 8'he5; ram[723] = 8'h21; 
    ram[724] = 8'h02; ram[725] = 8'h00; ram[726] = 8'h39; ram[727] = 8'hcd; 
    ram[728] = 8'h0d; ram[729] = 8'h00; ram[730] = 8'hd1; ram[731] = 8'h19; 
    ram[732] = 8'he5; ram[733] = 8'hcd; ram[734] = 8'h31; ram[735] = 8'h01; 
    ram[736] = 8'hc1; ram[737] = 8'hc1; ram[738] = 8'hc9; ram[739] = 8'h21; 
    ram[740] = 8'hc3; ram[741] = 8'h00; ram[742] = 8'h7d; ram[743] = 8'hd3; 
    ram[744] = 8'h81; ram[745] = 8'h21; ram[746] = 8'h00; ram[747] = 8'h00; 
    ram[748] = 8'h7d; ram[749] = 8'hd3; ram[750] = 8'h82; ram[751] = 8'h21; 
    ram[752] = 8'h5c; ram[753] = 8'h03; ram[754] = 8'he5; ram[755] = 8'hcd; 
    ram[756] = 8'h83; ram[757] = 8'h01; ram[758] = 8'hc1; ram[759] = 8'hcd; 
    ram[760] = 8'h72; ram[761] = 8'h01; ram[762] = 8'h21; ram[763] = 8'h6b; 
    ram[764] = 8'h03; ram[765] = 8'he5; ram[766] = 8'hcd; ram[767] = 8'h83; 
    ram[768] = 8'h01; ram[769] = 8'hc1; ram[770] = 8'h21; ram[771] = 8'h9f; 
    ram[772] = 8'h03; ram[773] = 8'he5; ram[774] = 8'h21; ram[775] = 8'h01; 
    ram[776] = 8'h00; ram[777] = 8'h29; ram[778] = 8'hd1; ram[779] = 8'h19; 
    ram[780] = 8'hcd; ram[781] = 8'h0d; ram[782] = 8'h00; ram[783] = 8'he5; 
    ram[784] = 8'hcd; ram[785] = 8'hb4; ram[786] = 8'h01; ram[787] = 8'hc1; 
    ram[788] = 8'hcd; ram[789] = 8'h72; ram[790] = 8'h01; ram[791] = 8'h21; 
    ram[792] = 8'h77; ram[793] = 8'h03; ram[794] = 8'he5; ram[795] = 8'hcd; 
    ram[796] = 8'h83; ram[797] = 8'h01; ram[798] = 8'hc1; ram[799] = 8'h21; 
    ram[800] = 8'h9f; ram[801] = 8'h03; ram[802] = 8'he5; ram[803] = 8'h21; 
    ram[804] = 8'h00; ram[805] = 8'h00; ram[806] = 8'h29; ram[807] = 8'hd1; 
    ram[808] = 8'h19; ram[809] = 8'hcd; ram[810] = 8'h0d; ram[811] = 8'h00; 
    ram[812] = 8'he5; ram[813] = 8'hcd; ram[814] = 8'h49; ram[815] = 8'h02; 
    ram[816] = 8'hc1; ram[817] = 8'hcd; ram[818] = 8'h72; ram[819] = 8'h01; 
    ram[820] = 8'h21; ram[821] = 8'h85; ram[822] = 8'h03; ram[823] = 8'he5; 
    ram[824] = 8'hcd; ram[825] = 8'h83; ram[826] = 8'h01; ram[827] = 8'hc1; 
    ram[828] = 8'hcd; ram[829] = 8'h72; ram[830] = 8'h01; ram[831] = 8'h21; 
    ram[832] = 8'h01; ram[833] = 8'h00; ram[834] = 8'h7c; ram[835] = 8'hb5; 
    ram[836] = 8'hca; ram[837] = 8'h5b; ram[838] = 8'h03; ram[839] = 8'hcd; 
    ram[840] = 8'h4f; ram[841] = 8'h01; ram[842] = 8'h7c; ram[843] = 8'hb5; 
    ram[844] = 8'hca; ram[845] = 8'h58; ram[846] = 8'h03; ram[847] = 8'h3a; 
    ram[848] = 8'h9e; ram[849] = 8'h03; ram[850] = 8'hcf; ram[851] = 8'he5; 
    ram[852] = 8'hcd; ram[853] = 8'h31; ram[854] = 8'h01; ram[855] = 8'hc1; 
    ram[856] = 8'hc3; ram[857] = 8'h3f; ram[858] = 8'h03; ram[859] = 8'hc9; 
    ram[860] = 8'h48; ram[861] = 8'h65; ram[862] = 8'h6c; ram[863] = 8'h6c; 
    ram[864] = 8'h6f; ram[865] = 8'h20; ram[866] = 8'h57; ram[867] = 8'h6f; 
    ram[868] = 8'h72; ram[869] = 8'h6c; ram[870] = 8'h64; ram[871] = 8'h21; 
    ram[872] = 8'h21; ram[873] = 8'h21; ram[874] = 8'h00; ram[875] = 8'h44; 
    ram[876] = 8'h65; ram[877] = 8'h63; ram[878] = 8'h20; ram[879] = 8'h76; 
    ram[880] = 8'h61; ram[881] = 8'h6c; ram[882] = 8'h75; ram[883] = 8'h65; 
    ram[884] = 8'h3a; ram[885] = 8'h20; ram[886] = 8'h00; ram[887] = 8'h48; 
    ram[888] = 8'h65; ram[889] = 8'h78; ram[890] = 8'h20; ram[891] = 8'h76; 
    ram[892] = 8'h61; ram[893] = 8'h6c; ram[894] = 8'h75; ram[895] = 8'h65; 
    ram[896] = 8'h3a; ram[897] = 8'h20; ram[898] = 8'h30; ram[899] = 8'h78; 
    ram[900] = 8'h00; ram[901] = 8'h45; ram[902] = 8'h63; ram[903] = 8'h68; 
    ram[904] = 8'h6f; ram[905] = 8'h69; ram[906] = 8'h6e; ram[907] = 8'h67; 
    ram[908] = 8'h20; ram[909] = 8'h72; ram[910] = 8'h65; ram[911] = 8'h63; 
    ram[912] = 8'h65; ram[913] = 8'h69; ram[914] = 8'h76; ram[915] = 8'h65; 
    ram[916] = 8'h64; ram[917] = 8'h20; ram[918] = 8'h62; ram[919] = 8'h79; 
    ram[920] = 8'h74; ram[921] = 8'h65; ram[922] = 8'h73; ram[923] = 8'h3a; 
    ram[924] = 8'h20; ram[925] = 8'h00; ram[926] = 8'h00; ram[927] = 8'hd2; 
    ram[928] = 8'h04; ram[929] = 8'h2e; ram[930] = 8'h16; ram[931] = 8'h00; 
    ram[932] = 8'h00; ram[933] = 8'h00; ram[934] = 8'h00; ram[935] = 8'h00; 
    ram[936] = 8'h00; ram[937] = 8'h00; ram[938] = 8'h00; ram[939] = 8'h00; 
    ram[940] = 8'h00; ram[941] = 8'h00; ram[942] = 8'h00; ram[943] = 8'h00; 
    ram[944] = 8'h00; ram[945] = 8'h00; ram[946] = 8'h00; ram[947] = 8'h00; 
    ram[948] = 8'h00; ram[949] = 8'h00; ram[950] = 8'h00; ram[951] = 8'h00; 
    ram[952] = 8'h00; ram[953] = 8'h00; ram[954] = 8'h00; ram[955] = 8'h00; 
    ram[956] = 8'h00; ram[957] = 8'h00; ram[958] = 8'h00; ram[959] = 8'h00; 
    ram[960] = 8'h00; ram[961] = 8'h00; ram[962] = 8'h00; ram[963] = 8'h00; 
    ram[964] = 8'h00; ram[965] = 8'h00; ram[966] = 8'h00; ram[967] = 8'h00; 
    ram[968] = 8'h00; ram[969] = 8'h00; ram[970] = 8'h00; ram[971] = 8'h00; 
    ram[972] = 8'h00; ram[973] = 8'h00; ram[974] = 8'h00; ram[975] = 8'h00; 
    ram[976] = 8'h00; ram[977] = 8'h00; ram[978] = 8'h00; ram[979] = 8'h00; 
    ram[980] = 8'h00; ram[981] = 8'h00; ram[982] = 8'h00; ram[983] = 8'h00; 
    ram[984] = 8'h00; ram[985] = 8'h00; ram[986] = 8'h00; ram[987] = 8'h00; 
    ram[988] = 8'h00; ram[989] = 8'h00; ram[990] = 8'h00; ram[991] = 8'h00; 
    ram[992] = 8'h00; ram[993] = 8'h00; ram[994] = 8'h00; ram[995] = 8'h00; 
    ram[996] = 8'h00; ram[997] = 8'h00; ram[998] = 8'h00; ram[999] = 8'h00; 
    ram[1000] = 8'h00; ram[1001] = 8'h00; ram[1002] = 8'h00; ram[1003] = 8'h00; 
    ram[1004] = 8'h00; ram[1005] = 8'h00; ram[1006] = 8'h00; ram[1007] = 8'h00; 
    ram[1008] = 8'h00; ram[1009] = 8'h00; ram[1010] = 8'h00; ram[1011] = 8'h00; 
    ram[1012] = 8'h00; ram[1013] = 8'h00; ram[1014] = 8'h00; ram[1015] = 8'h00; 
    ram[1016] = 8'h00; ram[1017] = 8'h00; ram[1018] = 8'h00; ram[1019] = 8'h00; 
    ram[1020] = 8'h00; ram[1021] = 8'h00; ram[1022] = 8'h00; ram[1023] = 8'h00; 
    ram[1024] = 8'h00; ram[1025] = 8'h00; ram[1026] = 8'h00; ram[1027] = 8'h00; 
    ram[1028] = 8'h00; ram[1029] = 8'h00; ram[1030] = 8'h00; ram[1031] = 8'h00; 
    ram[1032] = 8'h00; ram[1033] = 8'h00; ram[1034] = 8'h00; ram[1035] = 8'h00; 
    ram[1036] = 8'h00; ram[1037] = 8'h00; ram[1038] = 8'h00; ram[1039] = 8'h00; 
    ram[1040] = 8'h00; ram[1041] = 8'h00; ram[1042] = 8'h00; ram[1043] = 8'h00; 
    ram[1044] = 8'h00; ram[1045] = 8'h00; ram[1046] = 8'h00; ram[1047] = 8'h00; 
    ram[1048] = 8'h00; ram[1049] = 8'h00; ram[1050] = 8'h00; ram[1051] = 8'h00; 
    ram[1052] = 8'h00; ram[1053] = 8'h00; ram[1054] = 8'h00; ram[1055] = 8'h00; 
    ram[1056] = 8'h00; ram[1057] = 8'h00; ram[1058] = 8'h00; ram[1059] = 8'h00; 
    ram[1060] = 8'h00; ram[1061] = 8'h00; ram[1062] = 8'h00; ram[1063] = 8'h00; 
    ram[1064] = 8'h00; ram[1065] = 8'h00; ram[1066] = 8'h00; ram[1067] = 8'h00; 
    ram[1068] = 8'h00; ram[1069] = 8'h00; ram[1070] = 8'h00; ram[1071] = 8'h00; 
    ram[1072] = 8'h00; ram[1073] = 8'h00; ram[1074] = 8'h00; ram[1075] = 8'h00; 
    ram[1076] = 8'h00; ram[1077] = 8'h00; ram[1078] = 8'h00; ram[1079] = 8'h00; 
    ram[1080] = 8'h00; ram[1081] = 8'h00; ram[1082] = 8'h00; ram[1083] = 8'h00; 
    ram[1084] = 8'h00; ram[1085] = 8'h00; ram[1086] = 8'h00; ram[1087] = 8'h00; 
    ram[1088] = 8'h00; ram[1089] = 8'h00; ram[1090] = 8'h00; ram[1091] = 8'h00; 
    ram[1092] = 8'h00; ram[1093] = 8'h00; ram[1094] = 8'h00; ram[1095] = 8'h00; 
    ram[1096] = 8'h00; ram[1097] = 8'h00; ram[1098] = 8'h00; ram[1099] = 8'h00; 
    ram[1100] = 8'h00; ram[1101] = 8'h00; ram[1102] = 8'h00; ram[1103] = 8'h00; 
    ram[1104] = 8'h00; ram[1105] = 8'h00; ram[1106] = 8'h00; ram[1107] = 8'h00; 
    ram[1108] = 8'h00; ram[1109] = 8'h00; ram[1110] = 8'h00; ram[1111] = 8'h00; 
    ram[1112] = 8'h00; ram[1113] = 8'h00; ram[1114] = 8'h00; ram[1115] = 8'h00; 
    ram[1116] = 8'h00; ram[1117] = 8'h00; ram[1118] = 8'h00; ram[1119] = 8'h00; 
    ram[1120] = 8'h00; ram[1121] = 8'h00; ram[1122] = 8'h00; ram[1123] = 8'h00; 
    ram[1124] = 8'h00; ram[1125] = 8'h00; ram[1126] = 8'h00; ram[1127] = 8'h00; 
    ram[1128] = 8'h00; ram[1129] = 8'h00; ram[1130] = 8'h00; ram[1131] = 8'h00; 
    ram[1132] = 8'h00; ram[1133] = 8'h00; ram[1134] = 8'h00; ram[1135] = 8'h00; 
    ram[1136] = 8'h00; ram[1137] = 8'h00; ram[1138] = 8'h00; ram[1139] = 8'h00; 
    ram[1140] = 8'h00; ram[1141] = 8'h00; ram[1142] = 8'h00; ram[1143] = 8'h00; 
    ram[1144] = 8'h00; ram[1145] = 8'h00; ram[1146] = 8'h00; ram[1147] = 8'h00; 
    ram[1148] = 8'h00; ram[1149] = 8'h00; ram[1150] = 8'h00; ram[1151] = 8'h00; 
    ram[1152] = 8'h00; ram[1153] = 8'h00; ram[1154] = 8'h00; ram[1155] = 8'h00; 
    ram[1156] = 8'h00; ram[1157] = 8'h00; ram[1158] = 8'h00; ram[1159] = 8'h00; 
    ram[1160] = 8'h00; ram[1161] = 8'h00; ram[1162] = 8'h00; ram[1163] = 8'h00; 
    ram[1164] = 8'h00; ram[1165] = 8'h00; ram[1166] = 8'h00; ram[1167] = 8'h00; 
    ram[1168] = 8'h00; ram[1169] = 8'h00; ram[1170] = 8'h00; ram[1171] = 8'h00; 
    ram[1172] = 8'h00; ram[1173] = 8'h00; ram[1174] = 8'h00; ram[1175] = 8'h00; 
    ram[1176] = 8'h00; ram[1177] = 8'h00; ram[1178] = 8'h00; ram[1179] = 8'h00; 
    ram[1180] = 8'h00; ram[1181] = 8'h00; ram[1182] = 8'h00; ram[1183] = 8'h00; 
    ram[1184] = 8'h00; ram[1185] = 8'h00; ram[1186] = 8'h00; ram[1187] = 8'h00; 
    ram[1188] = 8'h00; ram[1189] = 8'h00; ram[1190] = 8'h00; ram[1191] = 8'h00; 
    ram[1192] = 8'h00; ram[1193] = 8'h00; ram[1194] = 8'h00; ram[1195] = 8'h00; 
    ram[1196] = 8'h00; ram[1197] = 8'h00; ram[1198] = 8'h00; ram[1199] = 8'h00; 
    ram[1200] = 8'h00; ram[1201] = 8'h00; ram[1202] = 8'h00; ram[1203] = 8'h00; 
    ram[1204] = 8'h00; ram[1205] = 8'h00; ram[1206] = 8'h00; ram[1207] = 8'h00; 
    ram[1208] = 8'h00; ram[1209] = 8'h00; ram[1210] = 8'h00; ram[1211] = 8'h00; 
    ram[1212] = 8'h00; ram[1213] = 8'h00; ram[1214] = 8'h00; ram[1215] = 8'h00; 
    ram[1216] = 8'h00; ram[1217] = 8'h00; ram[1218] = 8'h00; ram[1219] = 8'h00; 
    ram[1220] = 8'h00; ram[1221] = 8'h00; ram[1222] = 8'h00; ram[1223] = 8'h00; 
    ram[1224] = 8'h00; ram[1225] = 8'h00; ram[1226] = 8'h00; ram[1227] = 8'h00; 
    ram[1228] = 8'h00; ram[1229] = 8'h00; ram[1230] = 8'h00; ram[1231] = 8'h00; 
    ram[1232] = 8'h00; ram[1233] = 8'h00; ram[1234] = 8'h00; ram[1235] = 8'h00; 
    ram[1236] = 8'h00; ram[1237] = 8'h00; ram[1238] = 8'h00; ram[1239] = 8'h00; 
    ram[1240] = 8'h00; ram[1241] = 8'h00; ram[1242] = 8'h00; ram[1243] = 8'h00; 
    ram[1244] = 8'h00; ram[1245] = 8'h00; ram[1246] = 8'h00; ram[1247] = 8'h00; 
    ram[1248] = 8'h00; ram[1249] = 8'h00; ram[1250] = 8'h00; ram[1251] = 8'h00; 
    ram[1252] = 8'h00; ram[1253] = 8'h00; ram[1254] = 8'h00; ram[1255] = 8'h00; 
    ram[1256] = 8'h00; ram[1257] = 8'h00; ram[1258] = 8'h00; ram[1259] = 8'h00; 
    ram[1260] = 8'h00; ram[1261] = 8'h00; ram[1262] = 8'h00; ram[1263] = 8'h00; 
    ram[1264] = 8'h00; ram[1265] = 8'h00; ram[1266] = 8'h00; ram[1267] = 8'h00; 
    ram[1268] = 8'h00; ram[1269] = 8'h00; ram[1270] = 8'h00; ram[1271] = 8'h00; 
    ram[1272] = 8'h00; ram[1273] = 8'h00; ram[1274] = 8'h00; ram[1275] = 8'h00; 
    ram[1276] = 8'h00; ram[1277] = 8'h00; ram[1278] = 8'h00; ram[1279] = 8'h00; 
    ram[1280] = 8'h00; ram[1281] = 8'h00; ram[1282] = 8'h00; ram[1283] = 8'h00; 
    ram[1284] = 8'h00; ram[1285] = 8'h00; ram[1286] = 8'h00; ram[1287] = 8'h00; 
    ram[1288] = 8'h00; ram[1289] = 8'h00; ram[1290] = 8'h00; ram[1291] = 8'h00; 
    ram[1292] = 8'h00; ram[1293] = 8'h00; ram[1294] = 8'h00; ram[1295] = 8'h00; 
    ram[1296] = 8'h00; ram[1297] = 8'h00; ram[1298] = 8'h00; ram[1299] = 8'h00; 
    ram[1300] = 8'h00; ram[1301] = 8'h00; ram[1302] = 8'h00; ram[1303] = 8'h00; 
    ram[1304] = 8'h00; ram[1305] = 8'h00; ram[1306] = 8'h00; ram[1307] = 8'h00; 
    ram[1308] = 8'h00; ram[1309] = 8'h00; ram[1310] = 8'h00; ram[1311] = 8'h00; 
    ram[1312] = 8'h00; ram[1313] = 8'h00; ram[1314] = 8'h00; ram[1315] = 8'h00; 
    ram[1316] = 8'h00; ram[1317] = 8'h00; ram[1318] = 8'h00; ram[1319] = 8'h00; 
    ram[1320] = 8'h00; ram[1321] = 8'h00; ram[1322] = 8'h00; ram[1323] = 8'h00; 
    ram[1324] = 8'h00; ram[1325] = 8'h00; ram[1326] = 8'h00; ram[1327] = 8'h00; 
    ram[1328] = 8'h00; ram[1329] = 8'h00; ram[1330] = 8'h00; ram[1331] = 8'h00; 
    ram[1332] = 8'h00; ram[1333] = 8'h00; ram[1334] = 8'h00; ram[1335] = 8'h00; 
    ram[1336] = 8'h00; ram[1337] = 8'h00; ram[1338] = 8'h00; ram[1339] = 8'h00; 
    ram[1340] = 8'h00; ram[1341] = 8'h00; ram[1342] = 8'h00; ram[1343] = 8'h00; 
    ram[1344] = 8'h00; ram[1345] = 8'h00; ram[1346] = 8'h00; ram[1347] = 8'h00; 
    ram[1348] = 8'h00; ram[1349] = 8'h00; ram[1350] = 8'h00; ram[1351] = 8'h00; 
    ram[1352] = 8'h00; ram[1353] = 8'h00; ram[1354] = 8'h00; ram[1355] = 8'h00; 
    ram[1356] = 8'h00; ram[1357] = 8'h00; ram[1358] = 8'h00; ram[1359] = 8'h00; 
    ram[1360] = 8'h00; ram[1361] = 8'h00; ram[1362] = 8'h00; ram[1363] = 8'h00; 
    ram[1364] = 8'h00; ram[1365] = 8'h00; ram[1366] = 8'h00; ram[1367] = 8'h00; 
    ram[1368] = 8'h00; ram[1369] = 8'h00; ram[1370] = 8'h00; ram[1371] = 8'h00; 
    ram[1372] = 8'h00; ram[1373] = 8'h00; ram[1374] = 8'h00; ram[1375] = 8'h00; 
    ram[1376] = 8'h00; ram[1377] = 8'h00; ram[1378] = 8'h00; ram[1379] = 8'h00; 
    ram[1380] = 8'h00; ram[1381] = 8'h00; ram[1382] = 8'h00; ram[1383] = 8'h00; 
    ram[1384] = 8'h00; ram[1385] = 8'h00; ram[1386] = 8'h00; ram[1387] = 8'h00; 
    ram[1388] = 8'h00; ram[1389] = 8'h00; ram[1390] = 8'h00; ram[1391] = 8'h00; 
    ram[1392] = 8'h00; ram[1393] = 8'h00; ram[1394] = 8'h00; ram[1395] = 8'h00; 
    ram[1396] = 8'h00; ram[1397] = 8'h00; ram[1398] = 8'h00; ram[1399] = 8'h00; 
    ram[1400] = 8'h00; ram[1401] = 8'h00; ram[1402] = 8'h00; ram[1403] = 8'h00; 
    ram[1404] = 8'h00; ram[1405] = 8'h00; ram[1406] = 8'h00; ram[1407] = 8'h00; 
    ram[1408] = 8'h00; ram[1409] = 8'h00; ram[1410] = 8'h00; ram[1411] = 8'h00; 
    ram[1412] = 8'h00; ram[1413] = 8'h00; ram[1414] = 8'h00; ram[1415] = 8'h00; 
    ram[1416] = 8'h00; ram[1417] = 8'h00; ram[1418] = 8'h00; ram[1419] = 8'h00; 
    ram[1420] = 8'h00; ram[1421] = 8'h00; ram[1422] = 8'h00; ram[1423] = 8'h00; 
    ram[1424] = 8'h00; ram[1425] = 8'h00; ram[1426] = 8'h00; ram[1427] = 8'h00; 
    ram[1428] = 8'h00; ram[1429] = 8'h00; ram[1430] = 8'h00; ram[1431] = 8'h00; 
    ram[1432] = 8'h00; ram[1433] = 8'h00; ram[1434] = 8'h00; ram[1435] = 8'h00; 
    ram[1436] = 8'h00; ram[1437] = 8'h00; ram[1438] = 8'h00; ram[1439] = 8'h00; 
    ram[1440] = 8'h00; ram[1441] = 8'h00; ram[1442] = 8'h00; ram[1443] = 8'h00; 
    ram[1444] = 8'h00; ram[1445] = 8'h00; ram[1446] = 8'h00; ram[1447] = 8'h00; 
    ram[1448] = 8'h00; ram[1449] = 8'h00; ram[1450] = 8'h00; ram[1451] = 8'h00; 
    ram[1452] = 8'h00; ram[1453] = 8'h00; ram[1454] = 8'h00; ram[1455] = 8'h00; 
    ram[1456] = 8'h00; ram[1457] = 8'h00; ram[1458] = 8'h00; ram[1459] = 8'h00; 
    ram[1460] = 8'h00; ram[1461] = 8'h00; ram[1462] = 8'h00; ram[1463] = 8'h00; 
    ram[1464] = 8'h00; ram[1465] = 8'h00; ram[1466] = 8'h00; ram[1467] = 8'h00; 
    ram[1468] = 8'h00; ram[1469] = 8'h00; ram[1470] = 8'h00; ram[1471] = 8'h00; 
    ram[1472] = 8'h00; ram[1473] = 8'h00; ram[1474] = 8'h00; ram[1475] = 8'h00; 
    ram[1476] = 8'h00; ram[1477] = 8'h00; ram[1478] = 8'h00; ram[1479] = 8'h00; 
    ram[1480] = 8'h00; ram[1481] = 8'h00; ram[1482] = 8'h00; ram[1483] = 8'h00; 
    ram[1484] = 8'h00; ram[1485] = 8'h00; ram[1486] = 8'h00; ram[1487] = 8'h00; 
    ram[1488] = 8'h00; ram[1489] = 8'h00; ram[1490] = 8'h00; ram[1491] = 8'h00; 
    ram[1492] = 8'h00; ram[1493] = 8'h00; ram[1494] = 8'h00; ram[1495] = 8'h00; 
    ram[1496] = 8'h00; ram[1497] = 8'h00; ram[1498] = 8'h00; ram[1499] = 8'h00; 
    ram[1500] = 8'h00; ram[1501] = 8'h00; ram[1502] = 8'h00; ram[1503] = 8'h00; 
    ram[1504] = 8'h00; ram[1505] = 8'h00; ram[1506] = 8'h00; ram[1507] = 8'h00; 
    ram[1508] = 8'h00; ram[1509] = 8'h00; ram[1510] = 8'h00; ram[1511] = 8'h00; 
    ram[1512] = 8'h00; ram[1513] = 8'h00; ram[1514] = 8'h00; ram[1515] = 8'h00; 
    ram[1516] = 8'h00; ram[1517] = 8'h00; ram[1518] = 8'h00; ram[1519] = 8'h00; 
    ram[1520] = 8'h00; ram[1521] = 8'h00; ram[1522] = 8'h00; ram[1523] = 8'h00; 
    ram[1524] = 8'h00; ram[1525] = 8'h00; ram[1526] = 8'h00; ram[1527] = 8'h00; 
    ram[1528] = 8'h00; ram[1529] = 8'h00; ram[1530] = 8'h00; ram[1531] = 8'h00; 
    ram[1532] = 8'h00; ram[1533] = 8'h00; ram[1534] = 8'h00; ram[1535] = 8'h00; 
    ram[1536] = 8'h00; ram[1537] = 8'h00; ram[1538] = 8'h00; ram[1539] = 8'h00; 
    ram[1540] = 8'h00; ram[1541] = 8'h00; ram[1542] = 8'h00; ram[1543] = 8'h00; 
    ram[1544] = 8'h00; ram[1545] = 8'h00; ram[1546] = 8'h00; ram[1547] = 8'h00; 
    ram[1548] = 8'h00; ram[1549] = 8'h00; ram[1550] = 8'h00; ram[1551] = 8'h00; 
    ram[1552] = 8'h00; ram[1553] = 8'h00; ram[1554] = 8'h00; ram[1555] = 8'h00; 
    ram[1556] = 8'h00; ram[1557] = 8'h00; ram[1558] = 8'h00; ram[1559] = 8'h00; 
    ram[1560] = 8'h00; ram[1561] = 8'h00; ram[1562] = 8'h00; ram[1563] = 8'h00; 
    ram[1564] = 8'h00; ram[1565] = 8'h00; ram[1566] = 8'h00; ram[1567] = 8'h00; 
    ram[1568] = 8'h00; ram[1569] = 8'h00; ram[1570] = 8'h00; ram[1571] = 8'h00; 
    ram[1572] = 8'h00; ram[1573] = 8'h00; ram[1574] = 8'h00; ram[1575] = 8'h00; 
    ram[1576] = 8'h00; ram[1577] = 8'h00; ram[1578] = 8'h00; ram[1579] = 8'h00; 
    ram[1580] = 8'h00; ram[1581] = 8'h00; ram[1582] = 8'h00; ram[1583] = 8'h00; 
    ram[1584] = 8'h00; ram[1585] = 8'h00; ram[1586] = 8'h00; ram[1587] = 8'h00; 
    ram[1588] = 8'h00; ram[1589] = 8'h00; ram[1590] = 8'h00; ram[1591] = 8'h00; 
    ram[1592] = 8'h00; ram[1593] = 8'h00; ram[1594] = 8'h00; ram[1595] = 8'h00; 
    ram[1596] = 8'h00; ram[1597] = 8'h00; ram[1598] = 8'h00; ram[1599] = 8'h00; 
    ram[1600] = 8'h00; ram[1601] = 8'h00; ram[1602] = 8'h00; ram[1603] = 8'h00; 
    ram[1604] = 8'h00; ram[1605] = 8'h00; ram[1606] = 8'h00; ram[1607] = 8'h00; 
    ram[1608] = 8'h00; ram[1609] = 8'h00; ram[1610] = 8'h00; ram[1611] = 8'h00; 
    ram[1612] = 8'h00; ram[1613] = 8'h00; ram[1614] = 8'h00; ram[1615] = 8'h00; 
    ram[1616] = 8'h00; ram[1617] = 8'h00; ram[1618] = 8'h00; ram[1619] = 8'h00; 
    ram[1620] = 8'h00; ram[1621] = 8'h00; ram[1622] = 8'h00; ram[1623] = 8'h00; 
    ram[1624] = 8'h00; ram[1625] = 8'h00; ram[1626] = 8'h00; ram[1627] = 8'h00; 
    ram[1628] = 8'h00; ram[1629] = 8'h00; ram[1630] = 8'h00; ram[1631] = 8'h00; 
    ram[1632] = 8'h00; ram[1633] = 8'h00; ram[1634] = 8'h00; ram[1635] = 8'h00; 
    ram[1636] = 8'h00; ram[1637] = 8'h00; ram[1638] = 8'h00; ram[1639] = 8'h00; 
    ram[1640] = 8'h00; ram[1641] = 8'h00; ram[1642] = 8'h00; ram[1643] = 8'h00; 
    ram[1644] = 8'h00; ram[1645] = 8'h00; ram[1646] = 8'h00; ram[1647] = 8'h00; 
    ram[1648] = 8'h00; ram[1649] = 8'h00; ram[1650] = 8'h00; ram[1651] = 8'h00; 
    ram[1652] = 8'h00; ram[1653] = 8'h00; ram[1654] = 8'h00; ram[1655] = 8'h00; 
    ram[1656] = 8'h00; ram[1657] = 8'h00; ram[1658] = 8'h00; ram[1659] = 8'h00; 
    ram[1660] = 8'h00; ram[1661] = 8'h00; ram[1662] = 8'h00; ram[1663] = 8'h00; 
    ram[1664] = 8'h00; ram[1665] = 8'h00; ram[1666] = 8'h00; ram[1667] = 8'h00; 
    ram[1668] = 8'h00; ram[1669] = 8'h00; ram[1670] = 8'h00; ram[1671] = 8'h00; 
    ram[1672] = 8'h00; ram[1673] = 8'h00; ram[1674] = 8'h00; ram[1675] = 8'h00; 
    ram[1676] = 8'h00; ram[1677] = 8'h00; ram[1678] = 8'h00; ram[1679] = 8'h00; 
    ram[1680] = 8'h00; ram[1681] = 8'h00; ram[1682] = 8'h00; ram[1683] = 8'h00; 
    ram[1684] = 8'h00; ram[1685] = 8'h00; ram[1686] = 8'h00; ram[1687] = 8'h00; 
    ram[1688] = 8'h00; ram[1689] = 8'h00; ram[1690] = 8'h00; ram[1691] = 8'h00; 
    ram[1692] = 8'h00; ram[1693] = 8'h00; ram[1694] = 8'h00; ram[1695] = 8'h00; 
    ram[1696] = 8'h00; ram[1697] = 8'h00; ram[1698] = 8'h00; ram[1699] = 8'h00; 
    ram[1700] = 8'h00; ram[1701] = 8'h00; ram[1702] = 8'h00; ram[1703] = 8'h00; 
    ram[1704] = 8'h00; ram[1705] = 8'h00; ram[1706] = 8'h00; ram[1707] = 8'h00; 
    ram[1708] = 8'h00; ram[1709] = 8'h00; ram[1710] = 8'h00; ram[1711] = 8'h00; 
    ram[1712] = 8'h00; ram[1713] = 8'h00; ram[1714] = 8'h00; ram[1715] = 8'h00; 
    ram[1716] = 8'h00; ram[1717] = 8'h00; ram[1718] = 8'h00; ram[1719] = 8'h00; 
    ram[1720] = 8'h00; ram[1721] = 8'h00; ram[1722] = 8'h00; ram[1723] = 8'h00; 
    ram[1724] = 8'h00; ram[1725] = 8'h00; ram[1726] = 8'h00; ram[1727] = 8'h00; 
    ram[1728] = 8'h00; ram[1729] = 8'h00; ram[1730] = 8'h00; ram[1731] = 8'h00; 
    ram[1732] = 8'h00; ram[1733] = 8'h00; ram[1734] = 8'h00; ram[1735] = 8'h00; 
    ram[1736] = 8'h00; ram[1737] = 8'h00; ram[1738] = 8'h00; ram[1739] = 8'h00; 
    ram[1740] = 8'h00; ram[1741] = 8'h00; ram[1742] = 8'h00; ram[1743] = 8'h00; 
    ram[1744] = 8'h00; ram[1745] = 8'h00; ram[1746] = 8'h00; ram[1747] = 8'h00; 
    ram[1748] = 8'h00; ram[1749] = 8'h00; ram[1750] = 8'h00; ram[1751] = 8'h00; 
    ram[1752] = 8'h00; ram[1753] = 8'h00; ram[1754] = 8'h00; ram[1755] = 8'h00; 
    ram[1756] = 8'h00; ram[1757] = 8'h00; ram[1758] = 8'h00; ram[1759] = 8'h00; 
    ram[1760] = 8'h00; ram[1761] = 8'h00; ram[1762] = 8'h00; ram[1763] = 8'h00; 
    ram[1764] = 8'h00; ram[1765] = 8'h00; ram[1766] = 8'h00; ram[1767] = 8'h00; 
    ram[1768] = 8'h00; ram[1769] = 8'h00; ram[1770] = 8'h00; ram[1771] = 8'h00; 
    ram[1772] = 8'h00; ram[1773] = 8'h00; ram[1774] = 8'h00; ram[1775] = 8'h00; 
    ram[1776] = 8'h00; ram[1777] = 8'h00; ram[1778] = 8'h00; ram[1779] = 8'h00; 
    ram[1780] = 8'h00; ram[1781] = 8'h00; ram[1782] = 8'h00; ram[1783] = 8'h00; 
    ram[1784] = 8'h00; ram[1785] = 8'h00; ram[1786] = 8'h00; ram[1787] = 8'h00; 
    ram[1788] = 8'h00; ram[1789] = 8'h00; ram[1790] = 8'h00; ram[1791] = 8'h00; 
    ram[1792] = 8'h00; ram[1793] = 8'h00; ram[1794] = 8'h00; ram[1795] = 8'h00; 
    ram[1796] = 8'h00; ram[1797] = 8'h00; ram[1798] = 8'h00; ram[1799] = 8'h00; 
    ram[1800] = 8'h00; ram[1801] = 8'h00; ram[1802] = 8'h00; ram[1803] = 8'h00; 
    ram[1804] = 8'h00; ram[1805] = 8'h00; ram[1806] = 8'h00; ram[1807] = 8'h00; 
    ram[1808] = 8'h00; ram[1809] = 8'h00; ram[1810] = 8'h00; ram[1811] = 8'h00; 
    ram[1812] = 8'h00; ram[1813] = 8'h00; ram[1814] = 8'h00; ram[1815] = 8'h00; 
    ram[1816] = 8'h00; ram[1817] = 8'h00; ram[1818] = 8'h00; ram[1819] = 8'h00; 
    ram[1820] = 8'h00; ram[1821] = 8'h00; ram[1822] = 8'h00; ram[1823] = 8'h00; 
    ram[1824] = 8'h00; ram[1825] = 8'h00; ram[1826] = 8'h00; ram[1827] = 8'h00; 
    ram[1828] = 8'h00; ram[1829] = 8'h00; ram[1830] = 8'h00; ram[1831] = 8'h00; 
    ram[1832] = 8'h00; ram[1833] = 8'h00; ram[1834] = 8'h00; ram[1835] = 8'h00; 
    ram[1836] = 8'h00; ram[1837] = 8'h00; ram[1838] = 8'h00; ram[1839] = 8'h00; 
    ram[1840] = 8'h00; ram[1841] = 8'h00; ram[1842] = 8'h00; ram[1843] = 8'h00; 
    ram[1844] = 8'h00; ram[1845] = 8'h00; ram[1846] = 8'h00; ram[1847] = 8'h00; 
    ram[1848] = 8'h00; ram[1849] = 8'h00; ram[1850] = 8'h00; ram[1851] = 8'h00; 
    ram[1852] = 8'h00; ram[1853] = 8'h00; ram[1854] = 8'h00; ram[1855] = 8'h00; 
    ram[1856] = 8'h00; ram[1857] = 8'h00; ram[1858] = 8'h00; ram[1859] = 8'h00; 
    ram[1860] = 8'h00; ram[1861] = 8'h00; ram[1862] = 8'h00; ram[1863] = 8'h00; 
    ram[1864] = 8'h00; ram[1865] = 8'h00; ram[1866] = 8'h00; ram[1867] = 8'h00; 
    ram[1868] = 8'h00; ram[1869] = 8'h00; ram[1870] = 8'h00; ram[1871] = 8'h00; 
    ram[1872] = 8'h00; ram[1873] = 8'h00; ram[1874] = 8'h00; ram[1875] = 8'h00; 
    ram[1876] = 8'h00; ram[1877] = 8'h00; ram[1878] = 8'h00; ram[1879] = 8'h00; 
    ram[1880] = 8'h00; ram[1881] = 8'h00; ram[1882] = 8'h00; ram[1883] = 8'h00; 
    ram[1884] = 8'h00; ram[1885] = 8'h00; ram[1886] = 8'h00; ram[1887] = 8'h00; 
    ram[1888] = 8'h00; ram[1889] = 8'h00; ram[1890] = 8'h00; ram[1891] = 8'h00; 
    ram[1892] = 8'h00; ram[1893] = 8'h00; ram[1894] = 8'h00; ram[1895] = 8'h00; 
    ram[1896] = 8'h00; ram[1897] = 8'h00; ram[1898] = 8'h00; ram[1899] = 8'h00; 
    ram[1900] = 8'h00; ram[1901] = 8'h00; ram[1902] = 8'h00; ram[1903] = 8'h00; 
    ram[1904] = 8'h00; ram[1905] = 8'h00; ram[1906] = 8'h00; ram[1907] = 8'h00; 
    ram[1908] = 8'h00; ram[1909] = 8'h00; ram[1910] = 8'h00; ram[1911] = 8'h00; 
    ram[1912] = 8'h00; ram[1913] = 8'h00; ram[1914] = 8'h00; ram[1915] = 8'h00; 
    ram[1916] = 8'h00; ram[1917] = 8'h00; ram[1918] = 8'h00; ram[1919] = 8'h00; 
    ram[1920] = 8'h00; ram[1921] = 8'h00; ram[1922] = 8'h00; ram[1923] = 8'h00; 
    ram[1924] = 8'h00; ram[1925] = 8'h00; ram[1926] = 8'h00; ram[1927] = 8'h00; 
    ram[1928] = 8'h00; ram[1929] = 8'h00; ram[1930] = 8'h00; ram[1931] = 8'h00; 
    ram[1932] = 8'h00; ram[1933] = 8'h00; ram[1934] = 8'h00; ram[1935] = 8'h00; 
    ram[1936] = 8'h00; ram[1937] = 8'h00; ram[1938] = 8'h00; ram[1939] = 8'h00; 
    ram[1940] = 8'h00; ram[1941] = 8'h00; ram[1942] = 8'h00; ram[1943] = 8'h00; 
    ram[1944] = 8'h00; ram[1945] = 8'h00; ram[1946] = 8'h00; ram[1947] = 8'h00; 
    ram[1948] = 8'h00; ram[1949] = 8'h00; ram[1950] = 8'h00; ram[1951] = 8'h00; 
    ram[1952] = 8'h00; ram[1953] = 8'h00; ram[1954] = 8'h00; ram[1955] = 8'h00; 
    ram[1956] = 8'h00; ram[1957] = 8'h00; ram[1958] = 8'h00; ram[1959] = 8'h00; 
    ram[1960] = 8'h00; ram[1961] = 8'h00; ram[1962] = 8'h00; ram[1963] = 8'h00; 
    ram[1964] = 8'h00; ram[1965] = 8'h00; ram[1966] = 8'h00; ram[1967] = 8'h00; 
    ram[1968] = 8'h00; ram[1969] = 8'h00; ram[1970] = 8'h00; ram[1971] = 8'h00; 
    ram[1972] = 8'h00; ram[1973] = 8'h00; ram[1974] = 8'h00; ram[1975] = 8'h00; 
    ram[1976] = 8'h00; ram[1977] = 8'h00; ram[1978] = 8'h00; ram[1979] = 8'h00; 
    ram[1980] = 8'h00; ram[1981] = 8'h00; ram[1982] = 8'h00; ram[1983] = 8'h00; 
    ram[1984] = 8'h00; ram[1985] = 8'h00; ram[1986] = 8'h00; ram[1987] = 8'h00; 
    ram[1988] = 8'h00; ram[1989] = 8'h00; ram[1990] = 8'h00; ram[1991] = 8'h00; 
    ram[1992] = 8'h00; ram[1993] = 8'h00; ram[1994] = 8'h00; ram[1995] = 8'h00; 
    ram[1996] = 8'h00; ram[1997] = 8'h00; ram[1998] = 8'h00; ram[1999] = 8'h00; 
    ram[2000] = 8'h00; ram[2001] = 8'h00; ram[2002] = 8'h00; ram[2003] = 8'h00; 
    ram[2004] = 8'h00; ram[2005] = 8'h00; ram[2006] = 8'h00; ram[2007] = 8'h00; 
    ram[2008] = 8'h00; ram[2009] = 8'h00; ram[2010] = 8'h00; ram[2011] = 8'h00; 
    ram[2012] = 8'h00; ram[2013] = 8'h00; ram[2014] = 8'h00; ram[2015] = 8'h00; 
    ram[2016] = 8'h00; ram[2017] = 8'h00; ram[2018] = 8'h00; ram[2019] = 8'h00; 
    ram[2020] = 8'h00; ram[2021] = 8'h00; ram[2022] = 8'h00; ram[2023] = 8'h00; 
    ram[2024] = 8'h00; ram[2025] = 8'h00; ram[2026] = 8'h00; ram[2027] = 8'h00; 
    ram[2028] = 8'h00; ram[2029] = 8'h00; ram[2030] = 8'h00; ram[2031] = 8'h00; 
    ram[2032] = 8'h00; ram[2033] = 8'h00; ram[2034] = 8'h00; ram[2035] = 8'h00; 
    ram[2036] = 8'h00; ram[2037] = 8'h00; ram[2038] = 8'h00; ram[2039] = 8'h00; 
    ram[2040] = 8'h00; ram[2041] = 8'h00; ram[2042] = 8'h00; ram[2043] = 8'h00; 
    ram[2044] = 8'h00; ram[2045] = 8'h00; ram[2046] = 8'h00; ram[2047] = 8'h00; 
    ram[2048] = 8'h00; ram[2049] = 8'h00; ram[2050] = 8'h00; ram[2051] = 8'h00; 
    ram[2052] = 8'h00; ram[2053] = 8'h00; ram[2054] = 8'h00; ram[2055] = 8'h00; 
    ram[2056] = 8'h00; ram[2057] = 8'h00; ram[2058] = 8'h00; ram[2059] = 8'h00; 
    ram[2060] = 8'h00; ram[2061] = 8'h00; ram[2062] = 8'h00; ram[2063] = 8'h00; 
    ram[2064] = 8'h00; ram[2065] = 8'h00; ram[2066] = 8'h00; ram[2067] = 8'h00; 
    ram[2068] = 8'h00; ram[2069] = 8'h00; ram[2070] = 8'h00; ram[2071] = 8'h00; 
    ram[2072] = 8'h00; ram[2073] = 8'h00; ram[2074] = 8'h00; ram[2075] = 8'h00; 
    ram[2076] = 8'h00; ram[2077] = 8'h00; ram[2078] = 8'h00; ram[2079] = 8'h00; 
    ram[2080] = 8'h00; ram[2081] = 8'h00; ram[2082] = 8'h00; ram[2083] = 8'h00; 
    ram[2084] = 8'h00; ram[2085] = 8'h00; ram[2086] = 8'h00; ram[2087] = 8'h00; 
    ram[2088] = 8'h00; ram[2089] = 8'h00; ram[2090] = 8'h00; ram[2091] = 8'h00; 
    ram[2092] = 8'h00; ram[2093] = 8'h00; ram[2094] = 8'h00; ram[2095] = 8'h00; 
    ram[2096] = 8'h00; ram[2097] = 8'h00; ram[2098] = 8'h00; ram[2099] = 8'h00; 
    ram[2100] = 8'h00; ram[2101] = 8'h00; ram[2102] = 8'h00; ram[2103] = 8'h00; 
    ram[2104] = 8'h00; ram[2105] = 8'h00; ram[2106] = 8'h00; ram[2107] = 8'h00; 
    ram[2108] = 8'h00; ram[2109] = 8'h00; ram[2110] = 8'h00; ram[2111] = 8'h00; 
    ram[2112] = 8'h00; ram[2113] = 8'h00; ram[2114] = 8'h00; ram[2115] = 8'h00; 
    ram[2116] = 8'h00; ram[2117] = 8'h00; ram[2118] = 8'h00; ram[2119] = 8'h00; 
    ram[2120] = 8'h00; ram[2121] = 8'h00; ram[2122] = 8'h00; ram[2123] = 8'h00; 
    ram[2124] = 8'h00; ram[2125] = 8'h00; ram[2126] = 8'h00; ram[2127] = 8'h00; 
    ram[2128] = 8'h00; ram[2129] = 8'h00; ram[2130] = 8'h00; ram[2131] = 8'h00; 
    ram[2132] = 8'h00; ram[2133] = 8'h00; ram[2134] = 8'h00; ram[2135] = 8'h00; 
    ram[2136] = 8'h00; ram[2137] = 8'h00; ram[2138] = 8'h00; ram[2139] = 8'h00; 
    ram[2140] = 8'h00; ram[2141] = 8'h00; ram[2142] = 8'h00; ram[2143] = 8'h00; 
    ram[2144] = 8'h00; ram[2145] = 8'h00; ram[2146] = 8'h00; ram[2147] = 8'h00; 
    ram[2148] = 8'h00; ram[2149] = 8'h00; ram[2150] = 8'h00; ram[2151] = 8'h00; 
    ram[2152] = 8'h00; ram[2153] = 8'h00; ram[2154] = 8'h00; ram[2155] = 8'h00; 
    ram[2156] = 8'h00; ram[2157] = 8'h00; ram[2158] = 8'h00; ram[2159] = 8'h00; 
    ram[2160] = 8'h00; ram[2161] = 8'h00; ram[2162] = 8'h00; ram[2163] = 8'h00; 
    ram[2164] = 8'h00; ram[2165] = 8'h00; ram[2166] = 8'h00; ram[2167] = 8'h00; 
    ram[2168] = 8'h00; ram[2169] = 8'h00; ram[2170] = 8'h00; ram[2171] = 8'h00; 
    ram[2172] = 8'h00; ram[2173] = 8'h00; ram[2174] = 8'h00; ram[2175] = 8'h00; 
    ram[2176] = 8'h00; ram[2177] = 8'h00; ram[2178] = 8'h00; ram[2179] = 8'h00; 
    ram[2180] = 8'h00; ram[2181] = 8'h00; ram[2182] = 8'h00; ram[2183] = 8'h00; 
    ram[2184] = 8'h00; ram[2185] = 8'h00; ram[2186] = 8'h00; ram[2187] = 8'h00; 
    ram[2188] = 8'h00; ram[2189] = 8'h00; ram[2190] = 8'h00; ram[2191] = 8'h00; 
    ram[2192] = 8'h00; ram[2193] = 8'h00; ram[2194] = 8'h00; ram[2195] = 8'h00; 
    ram[2196] = 8'h00; ram[2197] = 8'h00; ram[2198] = 8'h00; ram[2199] = 8'h00; 
    ram[2200] = 8'h00; ram[2201] = 8'h00; ram[2202] = 8'h00; ram[2203] = 8'h00; 
    ram[2204] = 8'h00; ram[2205] = 8'h00; ram[2206] = 8'h00; ram[2207] = 8'h00; 
    ram[2208] = 8'h00; ram[2209] = 8'h00; ram[2210] = 8'h00; ram[2211] = 8'h00; 
    ram[2212] = 8'h00; ram[2213] = 8'h00; ram[2214] = 8'h00; ram[2215] = 8'h00; 
    ram[2216] = 8'h00; ram[2217] = 8'h00; ram[2218] = 8'h00; ram[2219] = 8'h00; 
    ram[2220] = 8'h00; ram[2221] = 8'h00; ram[2222] = 8'h00; ram[2223] = 8'h00; 
    ram[2224] = 8'h00; ram[2225] = 8'h00; ram[2226] = 8'h00; ram[2227] = 8'h00; 
    ram[2228] = 8'h00; ram[2229] = 8'h00; ram[2230] = 8'h00; ram[2231] = 8'h00; 
    ram[2232] = 8'h00; ram[2233] = 8'h00; ram[2234] = 8'h00; ram[2235] = 8'h00; 
    ram[2236] = 8'h00; ram[2237] = 8'h00; ram[2238] = 8'h00; ram[2239] = 8'h00; 
    ram[2240] = 8'h00; ram[2241] = 8'h00; ram[2242] = 8'h00; ram[2243] = 8'h00; 
    ram[2244] = 8'h00; ram[2245] = 8'h00; ram[2246] = 8'h00; ram[2247] = 8'h00; 
    ram[2248] = 8'h00; ram[2249] = 8'h00; ram[2250] = 8'h00; ram[2251] = 8'h00; 
    ram[2252] = 8'h00; ram[2253] = 8'h00; ram[2254] = 8'h00; ram[2255] = 8'h00; 
    ram[2256] = 8'h00; ram[2257] = 8'h00; ram[2258] = 8'h00; ram[2259] = 8'h00; 
    ram[2260] = 8'h00; ram[2261] = 8'h00; ram[2262] = 8'h00; ram[2263] = 8'h00; 
    ram[2264] = 8'h00; ram[2265] = 8'h00; ram[2266] = 8'h00; ram[2267] = 8'h00; 
    ram[2268] = 8'h00; ram[2269] = 8'h00; ram[2270] = 8'h00; ram[2271] = 8'h00; 
    ram[2272] = 8'h00; ram[2273] = 8'h00; ram[2274] = 8'h00; ram[2275] = 8'h00; 
    ram[2276] = 8'h00; ram[2277] = 8'h00; ram[2278] = 8'h00; ram[2279] = 8'h00; 
    ram[2280] = 8'h00; ram[2281] = 8'h00; ram[2282] = 8'h00; ram[2283] = 8'h00; 
    ram[2284] = 8'h00; ram[2285] = 8'h00; ram[2286] = 8'h00; ram[2287] = 8'h00; 
    ram[2288] = 8'h00; ram[2289] = 8'h00; ram[2290] = 8'h00; ram[2291] = 8'h00; 
    ram[2292] = 8'h00; ram[2293] = 8'h00; ram[2294] = 8'h00; ram[2295] = 8'h00; 
    ram[2296] = 8'h00; ram[2297] = 8'h00; ram[2298] = 8'h00; ram[2299] = 8'h00; 
    ram[2300] = 8'h00; ram[2301] = 8'h00; ram[2302] = 8'h00; ram[2303] = 8'h00; 
    ram[2304] = 8'h00; ram[2305] = 8'h00; ram[2306] = 8'h00; ram[2307] = 8'h00; 
    ram[2308] = 8'h00; ram[2309] = 8'h00; ram[2310] = 8'h00; ram[2311] = 8'h00; 
    ram[2312] = 8'h00; ram[2313] = 8'h00; ram[2314] = 8'h00; ram[2315] = 8'h00; 
    ram[2316] = 8'h00; ram[2317] = 8'h00; ram[2318] = 8'h00; ram[2319] = 8'h00; 
    ram[2320] = 8'h00; ram[2321] = 8'h00; ram[2322] = 8'h00; ram[2323] = 8'h00; 
    ram[2324] = 8'h00; ram[2325] = 8'h00; ram[2326] = 8'h00; ram[2327] = 8'h00; 
    ram[2328] = 8'h00; ram[2329] = 8'h00; ram[2330] = 8'h00; ram[2331] = 8'h00; 
    ram[2332] = 8'h00; ram[2333] = 8'h00; ram[2334] = 8'h00; ram[2335] = 8'h00; 
    ram[2336] = 8'h00; ram[2337] = 8'h00; ram[2338] = 8'h00; ram[2339] = 8'h00; 
    ram[2340] = 8'h00; ram[2341] = 8'h00; ram[2342] = 8'h00; ram[2343] = 8'h00; 
    ram[2344] = 8'h00; ram[2345] = 8'h00; ram[2346] = 8'h00; ram[2347] = 8'h00; 
    ram[2348] = 8'h00; ram[2349] = 8'h00; ram[2350] = 8'h00; ram[2351] = 8'h00; 
    ram[2352] = 8'h00; ram[2353] = 8'h00; ram[2354] = 8'h00; ram[2355] = 8'h00; 
    ram[2356] = 8'h00; ram[2357] = 8'h00; ram[2358] = 8'h00; ram[2359] = 8'h00; 
    ram[2360] = 8'h00; ram[2361] = 8'h00; ram[2362] = 8'h00; ram[2363] = 8'h00; 
    ram[2364] = 8'h00; ram[2365] = 8'h00; ram[2366] = 8'h00; ram[2367] = 8'h00; 
    ram[2368] = 8'h00; ram[2369] = 8'h00; ram[2370] = 8'h00; ram[2371] = 8'h00; 
    ram[2372] = 8'h00; ram[2373] = 8'h00; ram[2374] = 8'h00; ram[2375] = 8'h00; 
    ram[2376] = 8'h00; ram[2377] = 8'h00; ram[2378] = 8'h00; ram[2379] = 8'h00; 
    ram[2380] = 8'h00; ram[2381] = 8'h00; ram[2382] = 8'h00; ram[2383] = 8'h00; 
    ram[2384] = 8'h00; ram[2385] = 8'h00; ram[2386] = 8'h00; ram[2387] = 8'h00; 
    ram[2388] = 8'h00; ram[2389] = 8'h00; ram[2390] = 8'h00; ram[2391] = 8'h00; 
    ram[2392] = 8'h00; ram[2393] = 8'h00; ram[2394] = 8'h00; ram[2395] = 8'h00; 
    ram[2396] = 8'h00; ram[2397] = 8'h00; ram[2398] = 8'h00; ram[2399] = 8'h00; 
    ram[2400] = 8'h00; ram[2401] = 8'h00; ram[2402] = 8'h00; ram[2403] = 8'h00; 
    ram[2404] = 8'h00; ram[2405] = 8'h00; ram[2406] = 8'h00; ram[2407] = 8'h00; 
    ram[2408] = 8'h00; ram[2409] = 8'h00; ram[2410] = 8'h00; ram[2411] = 8'h00; 
    ram[2412] = 8'h00; ram[2413] = 8'h00; ram[2414] = 8'h00; ram[2415] = 8'h00; 
    ram[2416] = 8'h00; ram[2417] = 8'h00; ram[2418] = 8'h00; ram[2419] = 8'h00; 
    ram[2420] = 8'h00; ram[2421] = 8'h00; ram[2422] = 8'h00; ram[2423] = 8'h00; 
    ram[2424] = 8'h00; ram[2425] = 8'h00; ram[2426] = 8'h00; ram[2427] = 8'h00; 
    ram[2428] = 8'h00; ram[2429] = 8'h00; ram[2430] = 8'h00; ram[2431] = 8'h00; 
    ram[2432] = 8'h00; ram[2433] = 8'h00; ram[2434] = 8'h00; ram[2435] = 8'h00; 
    ram[2436] = 8'h00; ram[2437] = 8'h00; ram[2438] = 8'h00; ram[2439] = 8'h00; 
    ram[2440] = 8'h00; ram[2441] = 8'h00; ram[2442] = 8'h00; ram[2443] = 8'h00; 
    ram[2444] = 8'h00; ram[2445] = 8'h00; ram[2446] = 8'h00; ram[2447] = 8'h00; 
    ram[2448] = 8'h00; ram[2449] = 8'h00; ram[2450] = 8'h00; ram[2451] = 8'h00; 
    ram[2452] = 8'h00; ram[2453] = 8'h00; ram[2454] = 8'h00; ram[2455] = 8'h00; 
    ram[2456] = 8'h00; ram[2457] = 8'h00; ram[2458] = 8'h00; ram[2459] = 8'h00; 
    ram[2460] = 8'h00; ram[2461] = 8'h00; ram[2462] = 8'h00; ram[2463] = 8'h00; 
    ram[2464] = 8'h00; ram[2465] = 8'h00; ram[2466] = 8'h00; ram[2467] = 8'h00; 
    ram[2468] = 8'h00; ram[2469] = 8'h00; ram[2470] = 8'h00; ram[2471] = 8'h00; 
    ram[2472] = 8'h00; ram[2473] = 8'h00; ram[2474] = 8'h00; ram[2475] = 8'h00; 
    ram[2476] = 8'h00; ram[2477] = 8'h00; ram[2478] = 8'h00; ram[2479] = 8'h00; 
    ram[2480] = 8'h00; ram[2481] = 8'h00; ram[2482] = 8'h00; ram[2483] = 8'h00; 
    ram[2484] = 8'h00; ram[2485] = 8'h00; ram[2486] = 8'h00; ram[2487] = 8'h00; 
    ram[2488] = 8'h00; ram[2489] = 8'h00; ram[2490] = 8'h00; ram[2491] = 8'h00; 
    ram[2492] = 8'h00; ram[2493] = 8'h00; ram[2494] = 8'h00; ram[2495] = 8'h00; 
    ram[2496] = 8'h00; ram[2497] = 8'h00; ram[2498] = 8'h00; ram[2499] = 8'h00; 
    ram[2500] = 8'h00; ram[2501] = 8'h00; ram[2502] = 8'h00; ram[2503] = 8'h00; 
    ram[2504] = 8'h00; ram[2505] = 8'h00; ram[2506] = 8'h00; ram[2507] = 8'h00; 
    ram[2508] = 8'h00; ram[2509] = 8'h00; ram[2510] = 8'h00; ram[2511] = 8'h00; 
    ram[2512] = 8'h00; ram[2513] = 8'h00; ram[2514] = 8'h00; ram[2515] = 8'h00; 
    ram[2516] = 8'h00; ram[2517] = 8'h00; ram[2518] = 8'h00; ram[2519] = 8'h00; 
    ram[2520] = 8'h00; ram[2521] = 8'h00; ram[2522] = 8'h00; ram[2523] = 8'h00; 
    ram[2524] = 8'h00; ram[2525] = 8'h00; ram[2526] = 8'h00; ram[2527] = 8'h00; 
    ram[2528] = 8'h00; ram[2529] = 8'h00; ram[2530] = 8'h00; ram[2531] = 8'h00; 
    ram[2532] = 8'h00; ram[2533] = 8'h00; ram[2534] = 8'h00; ram[2535] = 8'h00; 
    ram[2536] = 8'h00; ram[2537] = 8'h00; ram[2538] = 8'h00; ram[2539] = 8'h00; 
    ram[2540] = 8'h00; ram[2541] = 8'h00; ram[2542] = 8'h00; ram[2543] = 8'h00; 
    ram[2544] = 8'h00; ram[2545] = 8'h00; ram[2546] = 8'h00; ram[2547] = 8'h00; 
    ram[2548] = 8'h00; ram[2549] = 8'h00; ram[2550] = 8'h00; ram[2551] = 8'h00; 
    ram[2552] = 8'h00; ram[2553] = 8'h00; ram[2554] = 8'h00; ram[2555] = 8'h00; 
    ram[2556] = 8'h00; ram[2557] = 8'h00; ram[2558] = 8'h00; ram[2559] = 8'h00; 
    ram[2560] = 8'h00; ram[2561] = 8'h00; ram[2562] = 8'h00; ram[2563] = 8'h00; 
    ram[2564] = 8'h00; ram[2565] = 8'h00; ram[2566] = 8'h00; ram[2567] = 8'h00; 
    ram[2568] = 8'h00; ram[2569] = 8'h00; ram[2570] = 8'h00; ram[2571] = 8'h00; 
    ram[2572] = 8'h00; ram[2573] = 8'h00; ram[2574] = 8'h00; ram[2575] = 8'h00; 
    ram[2576] = 8'h00; ram[2577] = 8'h00; ram[2578] = 8'h00; ram[2579] = 8'h00; 
    ram[2580] = 8'h00; ram[2581] = 8'h00; ram[2582] = 8'h00; ram[2583] = 8'h00; 
    ram[2584] = 8'h00; ram[2585] = 8'h00; ram[2586] = 8'h00; ram[2587] = 8'h00; 
    ram[2588] = 8'h00; ram[2589] = 8'h00; ram[2590] = 8'h00; ram[2591] = 8'h00; 
    ram[2592] = 8'h00; ram[2593] = 8'h00; ram[2594] = 8'h00; ram[2595] = 8'h00; 
    ram[2596] = 8'h00; ram[2597] = 8'h00; ram[2598] = 8'h00; ram[2599] = 8'h00; 
    ram[2600] = 8'h00; ram[2601] = 8'h00; ram[2602] = 8'h00; ram[2603] = 8'h00; 
    ram[2604] = 8'h00; ram[2605] = 8'h00; ram[2606] = 8'h00; ram[2607] = 8'h00; 
    ram[2608] = 8'h00; ram[2609] = 8'h00; ram[2610] = 8'h00; ram[2611] = 8'h00; 
    ram[2612] = 8'h00; ram[2613] = 8'h00; ram[2614] = 8'h00; ram[2615] = 8'h00; 
    ram[2616] = 8'h00; ram[2617] = 8'h00; ram[2618] = 8'h00; ram[2619] = 8'h00; 
    ram[2620] = 8'h00; ram[2621] = 8'h00; ram[2622] = 8'h00; ram[2623] = 8'h00; 
    ram[2624] = 8'h00; ram[2625] = 8'h00; ram[2626] = 8'h00; ram[2627] = 8'h00; 
    ram[2628] = 8'h00; ram[2629] = 8'h00; ram[2630] = 8'h00; ram[2631] = 8'h00; 
    ram[2632] = 8'h00; ram[2633] = 8'h00; ram[2634] = 8'h00; ram[2635] = 8'h00; 
    ram[2636] = 8'h00; ram[2637] = 8'h00; ram[2638] = 8'h00; ram[2639] = 8'h00; 
    ram[2640] = 8'h00; ram[2641] = 8'h00; ram[2642] = 8'h00; ram[2643] = 8'h00; 
    ram[2644] = 8'h00; ram[2645] = 8'h00; ram[2646] = 8'h00; ram[2647] = 8'h00; 
    ram[2648] = 8'h00; ram[2649] = 8'h00; ram[2650] = 8'h00; ram[2651] = 8'h00; 
    ram[2652] = 8'h00; ram[2653] = 8'h00; ram[2654] = 8'h00; ram[2655] = 8'h00; 
    ram[2656] = 8'h00; ram[2657] = 8'h00; ram[2658] = 8'h00; ram[2659] = 8'h00; 
    ram[2660] = 8'h00; ram[2661] = 8'h00; ram[2662] = 8'h00; ram[2663] = 8'h00; 
    ram[2664] = 8'h00; ram[2665] = 8'h00; ram[2666] = 8'h00; ram[2667] = 8'h00; 
    ram[2668] = 8'h00; ram[2669] = 8'h00; ram[2670] = 8'h00; ram[2671] = 8'h00; 
    ram[2672] = 8'h00; ram[2673] = 8'h00; ram[2674] = 8'h00; ram[2675] = 8'h00; 
    ram[2676] = 8'h00; ram[2677] = 8'h00; ram[2678] = 8'h00; ram[2679] = 8'h00; 
    ram[2680] = 8'h00; ram[2681] = 8'h00; ram[2682] = 8'h00; ram[2683] = 8'h00; 
    ram[2684] = 8'h00; ram[2685] = 8'h00; ram[2686] = 8'h00; ram[2687] = 8'h00; 
    ram[2688] = 8'h00; ram[2689] = 8'h00; ram[2690] = 8'h00; ram[2691] = 8'h00; 
    ram[2692] = 8'h00; ram[2693] = 8'h00; ram[2694] = 8'h00; ram[2695] = 8'h00; 
    ram[2696] = 8'h00; ram[2697] = 8'h00; ram[2698] = 8'h00; ram[2699] = 8'h00; 
    ram[2700] = 8'h00; ram[2701] = 8'h00; ram[2702] = 8'h00; ram[2703] = 8'h00; 
    ram[2704] = 8'h00; ram[2705] = 8'h00; ram[2706] = 8'h00; ram[2707] = 8'h00; 
    ram[2708] = 8'h00; ram[2709] = 8'h00; ram[2710] = 8'h00; ram[2711] = 8'h00; 
    ram[2712] = 8'h00; ram[2713] = 8'h00; ram[2714] = 8'h00; ram[2715] = 8'h00; 
    ram[2716] = 8'h00; ram[2717] = 8'h00; ram[2718] = 8'h00; ram[2719] = 8'h00; 
    ram[2720] = 8'h00; ram[2721] = 8'h00; ram[2722] = 8'h00; ram[2723] = 8'h00; 
    ram[2724] = 8'h00; ram[2725] = 8'h00; ram[2726] = 8'h00; ram[2727] = 8'h00; 
    ram[2728] = 8'h00; ram[2729] = 8'h00; ram[2730] = 8'h00; ram[2731] = 8'h00; 
    ram[2732] = 8'h00; ram[2733] = 8'h00; ram[2734] = 8'h00; ram[2735] = 8'h00; 
    ram[2736] = 8'h00; ram[2737] = 8'h00; ram[2738] = 8'h00; ram[2739] = 8'h00; 
    ram[2740] = 8'h00; ram[2741] = 8'h00; ram[2742] = 8'h00; ram[2743] = 8'h00; 
    ram[2744] = 8'h00; ram[2745] = 8'h00; ram[2746] = 8'h00; ram[2747] = 8'h00; 
    ram[2748] = 8'h00; ram[2749] = 8'h00; ram[2750] = 8'h00; ram[2751] = 8'h00; 
    ram[2752] = 8'h00; ram[2753] = 8'h00; ram[2754] = 8'h00; ram[2755] = 8'h00; 
    ram[2756] = 8'h00; ram[2757] = 8'h00; ram[2758] = 8'h00; ram[2759] = 8'h00; 
    ram[2760] = 8'h00; ram[2761] = 8'h00; ram[2762] = 8'h00; ram[2763] = 8'h00; 
    ram[2764] = 8'h00; ram[2765] = 8'h00; ram[2766] = 8'h00; ram[2767] = 8'h00; 
    ram[2768] = 8'h00; ram[2769] = 8'h00; ram[2770] = 8'h00; ram[2771] = 8'h00; 
    ram[2772] = 8'h00; ram[2773] = 8'h00; ram[2774] = 8'h00; ram[2775] = 8'h00; 
    ram[2776] = 8'h00; ram[2777] = 8'h00; ram[2778] = 8'h00; ram[2779] = 8'h00; 
    ram[2780] = 8'h00; ram[2781] = 8'h00; ram[2782] = 8'h00; ram[2783] = 8'h00; 
    ram[2784] = 8'h00; ram[2785] = 8'h00; ram[2786] = 8'h00; ram[2787] = 8'h00; 
    ram[2788] = 8'h00; ram[2789] = 8'h00; ram[2790] = 8'h00; ram[2791] = 8'h00; 
    ram[2792] = 8'h00; ram[2793] = 8'h00; ram[2794] = 8'h00; ram[2795] = 8'h00; 
    ram[2796] = 8'h00; ram[2797] = 8'h00; ram[2798] = 8'h00; ram[2799] = 8'h00; 
    ram[2800] = 8'h00; ram[2801] = 8'h00; ram[2802] = 8'h00; ram[2803] = 8'h00; 
    ram[2804] = 8'h00; ram[2805] = 8'h00; ram[2806] = 8'h00; ram[2807] = 8'h00; 
    ram[2808] = 8'h00; ram[2809] = 8'h00; ram[2810] = 8'h00; ram[2811] = 8'h00; 
    ram[2812] = 8'h00; ram[2813] = 8'h00; ram[2814] = 8'h00; ram[2815] = 8'h00; 
    ram[2816] = 8'h00; ram[2817] = 8'h00; ram[2818] = 8'h00; ram[2819] = 8'h00; 
    ram[2820] = 8'h00; ram[2821] = 8'h00; ram[2822] = 8'h00; ram[2823] = 8'h00; 
    ram[2824] = 8'h00; ram[2825] = 8'h00; ram[2826] = 8'h00; ram[2827] = 8'h00; 
    ram[2828] = 8'h00; ram[2829] = 8'h00; ram[2830] = 8'h00; ram[2831] = 8'h00; 
    ram[2832] = 8'h00; ram[2833] = 8'h00; ram[2834] = 8'h00; ram[2835] = 8'h00; 
    ram[2836] = 8'h00; ram[2837] = 8'h00; ram[2838] = 8'h00; ram[2839] = 8'h00; 
    ram[2840] = 8'h00; ram[2841] = 8'h00; ram[2842] = 8'h00; ram[2843] = 8'h00; 
    ram[2844] = 8'h00; ram[2845] = 8'h00; ram[2846] = 8'h00; ram[2847] = 8'h00; 
    ram[2848] = 8'h00; ram[2849] = 8'h00; ram[2850] = 8'h00; ram[2851] = 8'h00; 
    ram[2852] = 8'h00; ram[2853] = 8'h00; ram[2854] = 8'h00; ram[2855] = 8'h00; 
    ram[2856] = 8'h00; ram[2857] = 8'h00; ram[2858] = 8'h00; ram[2859] = 8'h00; 
    ram[2860] = 8'h00; ram[2861] = 8'h00; ram[2862] = 8'h00; ram[2863] = 8'h00; 
    ram[2864] = 8'h00; ram[2865] = 8'h00; ram[2866] = 8'h00; ram[2867] = 8'h00; 
    ram[2868] = 8'h00; ram[2869] = 8'h00; ram[2870] = 8'h00; ram[2871] = 8'h00; 
    ram[2872] = 8'h00; ram[2873] = 8'h00; ram[2874] = 8'h00; ram[2875] = 8'h00; 
    ram[2876] = 8'h00; ram[2877] = 8'h00; ram[2878] = 8'h00; ram[2879] = 8'h00; 
    ram[2880] = 8'h00; ram[2881] = 8'h00; ram[2882] = 8'h00; ram[2883] = 8'h00; 
    ram[2884] = 8'h00; ram[2885] = 8'h00; ram[2886] = 8'h00; ram[2887] = 8'h00; 
    ram[2888] = 8'h00; ram[2889] = 8'h00; ram[2890] = 8'h00; ram[2891] = 8'h00; 
    ram[2892] = 8'h00; ram[2893] = 8'h00; ram[2894] = 8'h00; ram[2895] = 8'h00; 
    ram[2896] = 8'h00; ram[2897] = 8'h00; ram[2898] = 8'h00; ram[2899] = 8'h00; 
    ram[2900] = 8'h00; ram[2901] = 8'h00; ram[2902] = 8'h00; ram[2903] = 8'h00; 
    ram[2904] = 8'h00; ram[2905] = 8'h00; ram[2906] = 8'h00; ram[2907] = 8'h00; 
    ram[2908] = 8'h00; ram[2909] = 8'h00; ram[2910] = 8'h00; ram[2911] = 8'h00; 
    ram[2912] = 8'h00; ram[2913] = 8'h00; ram[2914] = 8'h00; ram[2915] = 8'h00; 
    ram[2916] = 8'h00; ram[2917] = 8'h00; ram[2918] = 8'h00; ram[2919] = 8'h00; 
    ram[2920] = 8'h00; ram[2921] = 8'h00; ram[2922] = 8'h00; ram[2923] = 8'h00; 
    ram[2924] = 8'h00; ram[2925] = 8'h00; ram[2926] = 8'h00; ram[2927] = 8'h00; 
    ram[2928] = 8'h00; ram[2929] = 8'h00; ram[2930] = 8'h00; ram[2931] = 8'h00; 
    ram[2932] = 8'h00; ram[2933] = 8'h00; ram[2934] = 8'h00; ram[2935] = 8'h00; 
    ram[2936] = 8'h00; ram[2937] = 8'h00; ram[2938] = 8'h00; ram[2939] = 8'h00; 
    ram[2940] = 8'h00; ram[2941] = 8'h00; ram[2942] = 8'h00; ram[2943] = 8'h00; 
    ram[2944] = 8'h00; ram[2945] = 8'h00; ram[2946] = 8'h00; ram[2947] = 8'h00; 
    ram[2948] = 8'h00; ram[2949] = 8'h00; ram[2950] = 8'h00; ram[2951] = 8'h00; 
    ram[2952] = 8'h00; ram[2953] = 8'h00; ram[2954] = 8'h00; ram[2955] = 8'h00; 
    ram[2956] = 8'h00; ram[2957] = 8'h00; ram[2958] = 8'h00; ram[2959] = 8'h00; 
    ram[2960] = 8'h00; ram[2961] = 8'h00; ram[2962] = 8'h00; ram[2963] = 8'h00; 
    ram[2964] = 8'h00; ram[2965] = 8'h00; ram[2966] = 8'h00; ram[2967] = 8'h00; 
    ram[2968] = 8'h00; ram[2969] = 8'h00; ram[2970] = 8'h00; ram[2971] = 8'h00; 
    ram[2972] = 8'h00; ram[2973] = 8'h00; ram[2974] = 8'h00; ram[2975] = 8'h00; 
    ram[2976] = 8'h00; ram[2977] = 8'h00; ram[2978] = 8'h00; ram[2979] = 8'h00; 
    ram[2980] = 8'h00; ram[2981] = 8'h00; ram[2982] = 8'h00; ram[2983] = 8'h00; 
    ram[2984] = 8'h00; ram[2985] = 8'h00; ram[2986] = 8'h00; ram[2987] = 8'h00; 
    ram[2988] = 8'h00; ram[2989] = 8'h00; ram[2990] = 8'h00; ram[2991] = 8'h00; 
    ram[2992] = 8'h00; ram[2993] = 8'h00; ram[2994] = 8'h00; ram[2995] = 8'h00; 
    ram[2996] = 8'h00; ram[2997] = 8'h00; ram[2998] = 8'h00; ram[2999] = 8'h00; 
    ram[3000] = 8'h00; ram[3001] = 8'h00; ram[3002] = 8'h00; ram[3003] = 8'h00; 
    ram[3004] = 8'h00; ram[3005] = 8'h00; ram[3006] = 8'h00; ram[3007] = 8'h00; 
    ram[3008] = 8'h00; ram[3009] = 8'h00; ram[3010] = 8'h00; ram[3011] = 8'h00; 
    ram[3012] = 8'h00; ram[3013] = 8'h00; ram[3014] = 8'h00; ram[3015] = 8'h00; 
    ram[3016] = 8'h00; ram[3017] = 8'h00; ram[3018] = 8'h00; ram[3019] = 8'h00; 
    ram[3020] = 8'h00; ram[3021] = 8'h00; ram[3022] = 8'h00; ram[3023] = 8'h00; 
    ram[3024] = 8'h00; ram[3025] = 8'h00; ram[3026] = 8'h00; ram[3027] = 8'h00; 
    ram[3028] = 8'h00; ram[3029] = 8'h00; ram[3030] = 8'h00; ram[3031] = 8'h00; 
    ram[3032] = 8'h00; ram[3033] = 8'h00; ram[3034] = 8'h00; ram[3035] = 8'h00; 
    ram[3036] = 8'h00; ram[3037] = 8'h00; ram[3038] = 8'h00; ram[3039] = 8'h00; 
    ram[3040] = 8'h00; ram[3041] = 8'h00; ram[3042] = 8'h00; ram[3043] = 8'h00; 
    ram[3044] = 8'h00; ram[3045] = 8'h00; ram[3046] = 8'h00; ram[3047] = 8'h00; 
    ram[3048] = 8'h00; ram[3049] = 8'h00; ram[3050] = 8'h00; ram[3051] = 8'h00; 
    ram[3052] = 8'h00; ram[3053] = 8'h00; ram[3054] = 8'h00; ram[3055] = 8'h00; 
    ram[3056] = 8'h00; ram[3057] = 8'h00; ram[3058] = 8'h00; ram[3059] = 8'h00; 
    ram[3060] = 8'h00; ram[3061] = 8'h00; ram[3062] = 8'h00; ram[3063] = 8'h00; 
    ram[3064] = 8'h00; ram[3065] = 8'h00; ram[3066] = 8'h00; ram[3067] = 8'h00; 
    ram[3068] = 8'h00; ram[3069] = 8'h00; ram[3070] = 8'h00; ram[3071] = 8'h00; 
    ram[3072] = 8'h00; ram[3073] = 8'h00; ram[3074] = 8'h00; ram[3075] = 8'h00; 
    ram[3076] = 8'h00; ram[3077] = 8'h00; ram[3078] = 8'h00; ram[3079] = 8'h00; 
    ram[3080] = 8'h00; ram[3081] = 8'h00; ram[3082] = 8'h00; ram[3083] = 8'h00; 
    ram[3084] = 8'h00; ram[3085] = 8'h00; ram[3086] = 8'h00; ram[3087] = 8'h00; 
    ram[3088] = 8'h00; ram[3089] = 8'h00; ram[3090] = 8'h00; ram[3091] = 8'h00; 
    ram[3092] = 8'h00; ram[3093] = 8'h00; ram[3094] = 8'h00; ram[3095] = 8'h00; 
    ram[3096] = 8'h00; ram[3097] = 8'h00; ram[3098] = 8'h00; ram[3099] = 8'h00; 
    ram[3100] = 8'h00; ram[3101] = 8'h00; ram[3102] = 8'h00; ram[3103] = 8'h00; 
    ram[3104] = 8'h00; ram[3105] = 8'h00; ram[3106] = 8'h00; ram[3107] = 8'h00; 
    ram[3108] = 8'h00; ram[3109] = 8'h00; ram[3110] = 8'h00; ram[3111] = 8'h00; 
    ram[3112] = 8'h00; ram[3113] = 8'h00; ram[3114] = 8'h00; ram[3115] = 8'h00; 
    ram[3116] = 8'h00; ram[3117] = 8'h00; ram[3118] = 8'h00; ram[3119] = 8'h00; 
    ram[3120] = 8'h00; ram[3121] = 8'h00; ram[3122] = 8'h00; ram[3123] = 8'h00; 
    ram[3124] = 8'h00; ram[3125] = 8'h00; ram[3126] = 8'h00; ram[3127] = 8'h00; 
    ram[3128] = 8'h00; ram[3129] = 8'h00; ram[3130] = 8'h00; ram[3131] = 8'h00; 
    ram[3132] = 8'h00; ram[3133] = 8'h00; ram[3134] = 8'h00; ram[3135] = 8'h00; 
    ram[3136] = 8'h00; ram[3137] = 8'h00; ram[3138] = 8'h00; ram[3139] = 8'h00; 
    ram[3140] = 8'h00; ram[3141] = 8'h00; ram[3142] = 8'h00; ram[3143] = 8'h00; 
    ram[3144] = 8'h00; ram[3145] = 8'h00; ram[3146] = 8'h00; ram[3147] = 8'h00; 
    ram[3148] = 8'h00; ram[3149] = 8'h00; ram[3150] = 8'h00; ram[3151] = 8'h00; 
    ram[3152] = 8'h00; ram[3153] = 8'h00; ram[3154] = 8'h00; ram[3155] = 8'h00; 
    ram[3156] = 8'h00; ram[3157] = 8'h00; ram[3158] = 8'h00; ram[3159] = 8'h00; 
    ram[3160] = 8'h00; ram[3161] = 8'h00; ram[3162] = 8'h00; ram[3163] = 8'h00; 
    ram[3164] = 8'h00; ram[3165] = 8'h00; ram[3166] = 8'h00; ram[3167] = 8'h00; 
    ram[3168] = 8'h00; ram[3169] = 8'h00; ram[3170] = 8'h00; ram[3171] = 8'h00; 
    ram[3172] = 8'h00; ram[3173] = 8'h00; ram[3174] = 8'h00; ram[3175] = 8'h00; 
    ram[3176] = 8'h00; ram[3177] = 8'h00; ram[3178] = 8'h00; ram[3179] = 8'h00; 
    ram[3180] = 8'h00; ram[3181] = 8'h00; ram[3182] = 8'h00; ram[3183] = 8'h00; 
    ram[3184] = 8'h00; ram[3185] = 8'h00; ram[3186] = 8'h00; ram[3187] = 8'h00; 
    ram[3188] = 8'h00; ram[3189] = 8'h00; ram[3190] = 8'h00; ram[3191] = 8'h00; 
    ram[3192] = 8'h00; ram[3193] = 8'h00; ram[3194] = 8'h00; ram[3195] = 8'h00; 
    ram[3196] = 8'h00; ram[3197] = 8'h00; ram[3198] = 8'h00; ram[3199] = 8'h00; 
    ram[3200] = 8'h00; ram[3201] = 8'h00; ram[3202] = 8'h00; ram[3203] = 8'h00; 
    ram[3204] = 8'h00; ram[3205] = 8'h00; ram[3206] = 8'h00; ram[3207] = 8'h00; 
    ram[3208] = 8'h00; ram[3209] = 8'h00; ram[3210] = 8'h00; ram[3211] = 8'h00; 
    ram[3212] = 8'h00; ram[3213] = 8'h00; ram[3214] = 8'h00; ram[3215] = 8'h00; 
    ram[3216] = 8'h00; ram[3217] = 8'h00; ram[3218] = 8'h00; ram[3219] = 8'h00; 
    ram[3220] = 8'h00; ram[3221] = 8'h00; ram[3222] = 8'h00; ram[3223] = 8'h00; 
    ram[3224] = 8'h00; ram[3225] = 8'h00; ram[3226] = 8'h00; ram[3227] = 8'h00; 
    ram[3228] = 8'h00; ram[3229] = 8'h00; ram[3230] = 8'h00; ram[3231] = 8'h00; 
    ram[3232] = 8'h00; ram[3233] = 8'h00; ram[3234] = 8'h00; ram[3235] = 8'h00; 
    ram[3236] = 8'h00; ram[3237] = 8'h00; ram[3238] = 8'h00; ram[3239] = 8'h00; 
    ram[3240] = 8'h00; ram[3241] = 8'h00; ram[3242] = 8'h00; ram[3243] = 8'h00; 
    ram[3244] = 8'h00; ram[3245] = 8'h00; ram[3246] = 8'h00; ram[3247] = 8'h00; 
    ram[3248] = 8'h00; ram[3249] = 8'h00; ram[3250] = 8'h00; ram[3251] = 8'h00; 
    ram[3252] = 8'h00; ram[3253] = 8'h00; ram[3254] = 8'h00; ram[3255] = 8'h00; 
    ram[3256] = 8'h00; ram[3257] = 8'h00; ram[3258] = 8'h00; ram[3259] = 8'h00; 
    ram[3260] = 8'h00; ram[3261] = 8'h00; ram[3262] = 8'h00; ram[3263] = 8'h00; 
    ram[3264] = 8'h00; ram[3265] = 8'h00; ram[3266] = 8'h00; ram[3267] = 8'h00; 
    ram[3268] = 8'h00; ram[3269] = 8'h00; ram[3270] = 8'h00; ram[3271] = 8'h00; 
    ram[3272] = 8'h00; ram[3273] = 8'h00; ram[3274] = 8'h00; ram[3275] = 8'h00; 
    ram[3276] = 8'h00; ram[3277] = 8'h00; ram[3278] = 8'h00; ram[3279] = 8'h00; 
    ram[3280] = 8'h00; ram[3281] = 8'h00; ram[3282] = 8'h00; ram[3283] = 8'h00; 
    ram[3284] = 8'h00; ram[3285] = 8'h00; ram[3286] = 8'h00; ram[3287] = 8'h00; 
    ram[3288] = 8'h00; ram[3289] = 8'h00; ram[3290] = 8'h00; ram[3291] = 8'h00; 
    ram[3292] = 8'h00; ram[3293] = 8'h00; ram[3294] = 8'h00; ram[3295] = 8'h00; 
    ram[3296] = 8'h00; ram[3297] = 8'h00; ram[3298] = 8'h00; ram[3299] = 8'h00; 
    ram[3300] = 8'h00; ram[3301] = 8'h00; ram[3302] = 8'h00; ram[3303] = 8'h00; 
    ram[3304] = 8'h00; ram[3305] = 8'h00; ram[3306] = 8'h00; ram[3307] = 8'h00; 
    ram[3308] = 8'h00; ram[3309] = 8'h00; ram[3310] = 8'h00; ram[3311] = 8'h00; 
    ram[3312] = 8'h00; ram[3313] = 8'h00; ram[3314] = 8'h00; ram[3315] = 8'h00; 
    ram[3316] = 8'h00; ram[3317] = 8'h00; ram[3318] = 8'h00; ram[3319] = 8'h00; 
    ram[3320] = 8'h00; ram[3321] = 8'h00; ram[3322] = 8'h00; ram[3323] = 8'h00; 
    ram[3324] = 8'h00; ram[3325] = 8'h00; ram[3326] = 8'h00; ram[3327] = 8'h00; 
    ram[3328] = 8'h00; ram[3329] = 8'h00; ram[3330] = 8'h00; ram[3331] = 8'h00; 
    ram[3332] = 8'h00; ram[3333] = 8'h00; ram[3334] = 8'h00; ram[3335] = 8'h00; 
    ram[3336] = 8'h00; ram[3337] = 8'h00; ram[3338] = 8'h00; ram[3339] = 8'h00; 
    ram[3340] = 8'h00; ram[3341] = 8'h00; ram[3342] = 8'h00; ram[3343] = 8'h00; 
    ram[3344] = 8'h00; ram[3345] = 8'h00; ram[3346] = 8'h00; ram[3347] = 8'h00; 
    ram[3348] = 8'h00; ram[3349] = 8'h00; ram[3350] = 8'h00; ram[3351] = 8'h00; 
    ram[3352] = 8'h00; ram[3353] = 8'h00; ram[3354] = 8'h00; ram[3355] = 8'h00; 
    ram[3356] = 8'h00; ram[3357] = 8'h00; ram[3358] = 8'h00; ram[3359] = 8'h00; 
    ram[3360] = 8'h00; ram[3361] = 8'h00; ram[3362] = 8'h00; ram[3363] = 8'h00; 
    ram[3364] = 8'h00; ram[3365] = 8'h00; ram[3366] = 8'h00; ram[3367] = 8'h00; 
    ram[3368] = 8'h00; ram[3369] = 8'h00; ram[3370] = 8'h00; ram[3371] = 8'h00; 
    ram[3372] = 8'h00; ram[3373] = 8'h00; ram[3374] = 8'h00; ram[3375] = 8'h00; 
    ram[3376] = 8'h00; ram[3377] = 8'h00; ram[3378] = 8'h00; ram[3379] = 8'h00; 
    ram[3380] = 8'h00; ram[3381] = 8'h00; ram[3382] = 8'h00; ram[3383] = 8'h00; 
    ram[3384] = 8'h00; ram[3385] = 8'h00; ram[3386] = 8'h00; ram[3387] = 8'h00; 
    ram[3388] = 8'h00; ram[3389] = 8'h00; ram[3390] = 8'h00; ram[3391] = 8'h00; 
    ram[3392] = 8'h00; ram[3393] = 8'h00; ram[3394] = 8'h00; ram[3395] = 8'h00; 
    ram[3396] = 8'h00; ram[3397] = 8'h00; ram[3398] = 8'h00; ram[3399] = 8'h00; 
    ram[3400] = 8'h00; ram[3401] = 8'h00; ram[3402] = 8'h00; ram[3403] = 8'h00; 
    ram[3404] = 8'h00; ram[3405] = 8'h00; ram[3406] = 8'h00; ram[3407] = 8'h00; 
    ram[3408] = 8'h00; ram[3409] = 8'h00; ram[3410] = 8'h00; ram[3411] = 8'h00; 
    ram[3412] = 8'h00; ram[3413] = 8'h00; ram[3414] = 8'h00; ram[3415] = 8'h00; 
    ram[3416] = 8'h00; ram[3417] = 8'h00; ram[3418] = 8'h00; ram[3419] = 8'h00; 
    ram[3420] = 8'h00; ram[3421] = 8'h00; ram[3422] = 8'h00; ram[3423] = 8'h00; 
    ram[3424] = 8'h00; ram[3425] = 8'h00; ram[3426] = 8'h00; ram[3427] = 8'h00; 
    ram[3428] = 8'h00; ram[3429] = 8'h00; ram[3430] = 8'h00; ram[3431] = 8'h00; 
    ram[3432] = 8'h00; ram[3433] = 8'h00; ram[3434] = 8'h00; ram[3435] = 8'h00; 
    ram[3436] = 8'h00; ram[3437] = 8'h00; ram[3438] = 8'h00; ram[3439] = 8'h00; 
    ram[3440] = 8'h00; ram[3441] = 8'h00; ram[3442] = 8'h00; ram[3443] = 8'h00; 
    ram[3444] = 8'h00; ram[3445] = 8'h00; ram[3446] = 8'h00; ram[3447] = 8'h00; 
    ram[3448] = 8'h00; ram[3449] = 8'h00; ram[3450] = 8'h00; ram[3451] = 8'h00; 
    ram[3452] = 8'h00; ram[3453] = 8'h00; ram[3454] = 8'h00; ram[3455] = 8'h00; 
    ram[3456] = 8'h00; ram[3457] = 8'h00; ram[3458] = 8'h00; ram[3459] = 8'h00; 
    ram[3460] = 8'h00; ram[3461] = 8'h00; ram[3462] = 8'h00; ram[3463] = 8'h00; 
    ram[3464] = 8'h00; ram[3465] = 8'h00; ram[3466] = 8'h00; ram[3467] = 8'h00; 
    ram[3468] = 8'h00; ram[3469] = 8'h00; ram[3470] = 8'h00; ram[3471] = 8'h00; 
    ram[3472] = 8'h00; ram[3473] = 8'h00; ram[3474] = 8'h00; ram[3475] = 8'h00; 
    ram[3476] = 8'h00; ram[3477] = 8'h00; ram[3478] = 8'h00; ram[3479] = 8'h00; 
    ram[3480] = 8'h00; ram[3481] = 8'h00; ram[3482] = 8'h00; ram[3483] = 8'h00; 
    ram[3484] = 8'h00; ram[3485] = 8'h00; ram[3486] = 8'h00; ram[3487] = 8'h00; 
    ram[3488] = 8'h00; ram[3489] = 8'h00; ram[3490] = 8'h00; ram[3491] = 8'h00; 
    ram[3492] = 8'h00; ram[3493] = 8'h00; ram[3494] = 8'h00; ram[3495] = 8'h00; 
    ram[3496] = 8'h00; ram[3497] = 8'h00; ram[3498] = 8'h00; ram[3499] = 8'h00; 
    ram[3500] = 8'h00; ram[3501] = 8'h00; ram[3502] = 8'h00; ram[3503] = 8'h00; 
    ram[3504] = 8'h00; ram[3505] = 8'h00; ram[3506] = 8'h00; ram[3507] = 8'h00; 
    ram[3508] = 8'h00; ram[3509] = 8'h00; ram[3510] = 8'h00; ram[3511] = 8'h00; 
    ram[3512] = 8'h00; ram[3513] = 8'h00; ram[3514] = 8'h00; ram[3515] = 8'h00; 
    ram[3516] = 8'h00; ram[3517] = 8'h00; ram[3518] = 8'h00; ram[3519] = 8'h00; 
    ram[3520] = 8'h00; ram[3521] = 8'h00; ram[3522] = 8'h00; ram[3523] = 8'h00; 
    ram[3524] = 8'h00; ram[3525] = 8'h00; ram[3526] = 8'h00; ram[3527] = 8'h00; 
    ram[3528] = 8'h00; ram[3529] = 8'h00; ram[3530] = 8'h00; ram[3531] = 8'h00; 
    ram[3532] = 8'h00; ram[3533] = 8'h00; ram[3534] = 8'h00; ram[3535] = 8'h00; 
    ram[3536] = 8'h00; ram[3537] = 8'h00; ram[3538] = 8'h00; ram[3539] = 8'h00; 
    ram[3540] = 8'h00; ram[3541] = 8'h00; ram[3542] = 8'h00; ram[3543] = 8'h00; 
    ram[3544] = 8'h00; ram[3545] = 8'h00; ram[3546] = 8'h00; ram[3547] = 8'h00; 
    ram[3548] = 8'h00; ram[3549] = 8'h00; ram[3550] = 8'h00; ram[3551] = 8'h00; 
    ram[3552] = 8'h00; ram[3553] = 8'h00; ram[3554] = 8'h00; ram[3555] = 8'h00; 
    ram[3556] = 8'h00; ram[3557] = 8'h00; ram[3558] = 8'h00; ram[3559] = 8'h00; 
    ram[3560] = 8'h00; ram[3561] = 8'h00; ram[3562] = 8'h00; ram[3563] = 8'h00; 
    ram[3564] = 8'h00; ram[3565] = 8'h00; ram[3566] = 8'h00; ram[3567] = 8'h00; 
    ram[3568] = 8'h00; ram[3569] = 8'h00; ram[3570] = 8'h00; ram[3571] = 8'h00; 
    ram[3572] = 8'h00; ram[3573] = 8'h00; ram[3574] = 8'h00; ram[3575] = 8'h00; 
    ram[3576] = 8'h00; ram[3577] = 8'h00; ram[3578] = 8'h00; ram[3579] = 8'h00; 
    ram[3580] = 8'h00; ram[3581] = 8'h00; ram[3582] = 8'h00; ram[3583] = 8'h00; 
    ram[3584] = 8'h00; ram[3585] = 8'h00; ram[3586] = 8'h00; ram[3587] = 8'h00; 
    ram[3588] = 8'h00; ram[3589] = 8'h00; ram[3590] = 8'h00; ram[3591] = 8'h00; 
    ram[3592] = 8'h00; ram[3593] = 8'h00; ram[3594] = 8'h00; ram[3595] = 8'h00; 
    ram[3596] = 8'h00; ram[3597] = 8'h00; ram[3598] = 8'h00; ram[3599] = 8'h00; 
    ram[3600] = 8'h00; ram[3601] = 8'h00; ram[3602] = 8'h00; ram[3603] = 8'h00; 
    ram[3604] = 8'h00; ram[3605] = 8'h00; ram[3606] = 8'h00; ram[3607] = 8'h00; 
    ram[3608] = 8'h00; ram[3609] = 8'h00; ram[3610] = 8'h00; ram[3611] = 8'h00; 
    ram[3612] = 8'h00; ram[3613] = 8'h00; ram[3614] = 8'h00; ram[3615] = 8'h00; 
    ram[3616] = 8'h00; ram[3617] = 8'h00; ram[3618] = 8'h00; ram[3619] = 8'h00; 
    ram[3620] = 8'h00; ram[3621] = 8'h00; ram[3622] = 8'h00; ram[3623] = 8'h00; 
    ram[3624] = 8'h00; ram[3625] = 8'h00; ram[3626] = 8'h00; ram[3627] = 8'h00; 
    ram[3628] = 8'h00; ram[3629] = 8'h00; ram[3630] = 8'h00; ram[3631] = 8'h00; 
    ram[3632] = 8'h00; ram[3633] = 8'h00; ram[3634] = 8'h00; ram[3635] = 8'h00; 
    ram[3636] = 8'h00; ram[3637] = 8'h00; ram[3638] = 8'h00; ram[3639] = 8'h00; 
    ram[3640] = 8'h00; ram[3641] = 8'h00; ram[3642] = 8'h00; ram[3643] = 8'h00; 
    ram[3644] = 8'h00; ram[3645] = 8'h00; ram[3646] = 8'h00; ram[3647] = 8'h00; 
    ram[3648] = 8'h00; ram[3649] = 8'h00; ram[3650] = 8'h00; ram[3651] = 8'h00; 
    ram[3652] = 8'h00; ram[3653] = 8'h00; ram[3654] = 8'h00; ram[3655] = 8'h00; 
    ram[3656] = 8'h00; ram[3657] = 8'h00; ram[3658] = 8'h00; ram[3659] = 8'h00; 
    ram[3660] = 8'h00; ram[3661] = 8'h00; ram[3662] = 8'h00; ram[3663] = 8'h00; 
    ram[3664] = 8'h00; ram[3665] = 8'h00; ram[3666] = 8'h00; ram[3667] = 8'h00; 
    ram[3668] = 8'h00; ram[3669] = 8'h00; ram[3670] = 8'h00; ram[3671] = 8'h00; 
    ram[3672] = 8'h00; ram[3673] = 8'h00; ram[3674] = 8'h00; ram[3675] = 8'h00; 
    ram[3676] = 8'h00; ram[3677] = 8'h00; ram[3678] = 8'h00; ram[3679] = 8'h00; 
    ram[3680] = 8'h00; ram[3681] = 8'h00; ram[3682] = 8'h00; ram[3683] = 8'h00; 
    ram[3684] = 8'h00; ram[3685] = 8'h00; ram[3686] = 8'h00; ram[3687] = 8'h00; 
    ram[3688] = 8'h00; ram[3689] = 8'h00; ram[3690] = 8'h00; ram[3691] = 8'h00; 
    ram[3692] = 8'h00; ram[3693] = 8'h00; ram[3694] = 8'h00; ram[3695] = 8'h00; 
    ram[3696] = 8'h00; ram[3697] = 8'h00; ram[3698] = 8'h00; ram[3699] = 8'h00; 
    ram[3700] = 8'h00; ram[3701] = 8'h00; ram[3702] = 8'h00; ram[3703] = 8'h00; 
    ram[3704] = 8'h00; ram[3705] = 8'h00; ram[3706] = 8'h00; ram[3707] = 8'h00; 
    ram[3708] = 8'h00; ram[3709] = 8'h00; ram[3710] = 8'h00; ram[3711] = 8'h00; 
    ram[3712] = 8'h00; ram[3713] = 8'h00; ram[3714] = 8'h00; ram[3715] = 8'h00; 
    ram[3716] = 8'h00; ram[3717] = 8'h00; ram[3718] = 8'h00; ram[3719] = 8'h00; 
    ram[3720] = 8'h00; ram[3721] = 8'h00; ram[3722] = 8'h00; ram[3723] = 8'h00; 
    ram[3724] = 8'h00; ram[3725] = 8'h00; ram[3726] = 8'h00; ram[3727] = 8'h00; 
    ram[3728] = 8'h00; ram[3729] = 8'h00; ram[3730] = 8'h00; ram[3731] = 8'h00; 
    ram[3732] = 8'h00; ram[3733] = 8'h00; ram[3734] = 8'h00; ram[3735] = 8'h00; 
    ram[3736] = 8'h00; ram[3737] = 8'h00; ram[3738] = 8'h00; ram[3739] = 8'h00; 
    ram[3740] = 8'h00; ram[3741] = 8'h00; ram[3742] = 8'h00; ram[3743] = 8'h00; 
    ram[3744] = 8'h00; ram[3745] = 8'h00; ram[3746] = 8'h00; ram[3747] = 8'h00; 
    ram[3748] = 8'h00; ram[3749] = 8'h00; ram[3750] = 8'h00; ram[3751] = 8'h00; 
    ram[3752] = 8'h00; ram[3753] = 8'h00; ram[3754] = 8'h00; ram[3755] = 8'h00; 
    ram[3756] = 8'h00; ram[3757] = 8'h00; ram[3758] = 8'h00; ram[3759] = 8'h00; 
    ram[3760] = 8'h00; ram[3761] = 8'h00; ram[3762] = 8'h00; ram[3763] = 8'h00; 
    ram[3764] = 8'h00; ram[3765] = 8'h00; ram[3766] = 8'h00; ram[3767] = 8'h00; 
    ram[3768] = 8'h00; ram[3769] = 8'h00; ram[3770] = 8'h00; ram[3771] = 8'h00; 
    ram[3772] = 8'h00; ram[3773] = 8'h00; ram[3774] = 8'h00; ram[3775] = 8'h00; 
    ram[3776] = 8'h00; ram[3777] = 8'h00; ram[3778] = 8'h00; ram[3779] = 8'h00; 
    ram[3780] = 8'h00; ram[3781] = 8'h00; ram[3782] = 8'h00; ram[3783] = 8'h00; 
    ram[3784] = 8'h00; ram[3785] = 8'h00; ram[3786] = 8'h00; ram[3787] = 8'h00; 
    ram[3788] = 8'h00; ram[3789] = 8'h00; ram[3790] = 8'h00; ram[3791] = 8'h00; 
    ram[3792] = 8'h00; ram[3793] = 8'h00; ram[3794] = 8'h00; ram[3795] = 8'h00; 
    ram[3796] = 8'h00; ram[3797] = 8'h00; ram[3798] = 8'h00; ram[3799] = 8'h00; 
    ram[3800] = 8'h00; ram[3801] = 8'h00; ram[3802] = 8'h00; ram[3803] = 8'h00; 
    ram[3804] = 8'h00; ram[3805] = 8'h00; ram[3806] = 8'h00; ram[3807] = 8'h00; 
    ram[3808] = 8'h00; ram[3809] = 8'h00; ram[3810] = 8'h00; ram[3811] = 8'h00; 
    ram[3812] = 8'h00; ram[3813] = 8'h00; ram[3814] = 8'h00; ram[3815] = 8'h00; 
    ram[3816] = 8'h00; ram[3817] = 8'h00; ram[3818] = 8'h00; ram[3819] = 8'h00; 
    ram[3820] = 8'h00; ram[3821] = 8'h00; ram[3822] = 8'h00; ram[3823] = 8'h00; 
    ram[3824] = 8'h00; ram[3825] = 8'h00; ram[3826] = 8'h00; ram[3827] = 8'h00; 
    ram[3828] = 8'h00; ram[3829] = 8'h00; ram[3830] = 8'h00; ram[3831] = 8'h00; 
    ram[3832] = 8'h00; ram[3833] = 8'h00; ram[3834] = 8'h00; ram[3835] = 8'h00; 
    ram[3836] = 8'h00; ram[3837] = 8'h00; ram[3838] = 8'h00; ram[3839] = 8'h00; 
    ram[3840] = 8'h00; ram[3841] = 8'h00; ram[3842] = 8'h00; ram[3843] = 8'h00; 
    ram[3844] = 8'h00; ram[3845] = 8'h00; ram[3846] = 8'h00; ram[3847] = 8'h00; 
    ram[3848] = 8'h00; ram[3849] = 8'h00; ram[3850] = 8'h00; ram[3851] = 8'h00; 
    ram[3852] = 8'h00; ram[3853] = 8'h00; ram[3854] = 8'h00; ram[3855] = 8'h00; 
    ram[3856] = 8'h00; ram[3857] = 8'h00; ram[3858] = 8'h00; ram[3859] = 8'h00; 
    ram[3860] = 8'h00; ram[3861] = 8'h00; ram[3862] = 8'h00; ram[3863] = 8'h00; 
    ram[3864] = 8'h00; ram[3865] = 8'h00; ram[3866] = 8'h00; ram[3867] = 8'h00; 
    ram[3868] = 8'h00; ram[3869] = 8'h00; ram[3870] = 8'h00; ram[3871] = 8'h00; 
    ram[3872] = 8'h00; ram[3873] = 8'h00; ram[3874] = 8'h00; ram[3875] = 8'h00; 
    ram[3876] = 8'h00; ram[3877] = 8'h00; ram[3878] = 8'h00; ram[3879] = 8'h00; 
    ram[3880] = 8'h00; ram[3881] = 8'h00; ram[3882] = 8'h00; ram[3883] = 8'h00; 
    ram[3884] = 8'h00; ram[3885] = 8'h00; ram[3886] = 8'h00; ram[3887] = 8'h00; 
    ram[3888] = 8'h00; ram[3889] = 8'h00; ram[3890] = 8'h00; ram[3891] = 8'h00; 
    ram[3892] = 8'h00; ram[3893] = 8'h00; ram[3894] = 8'h00; ram[3895] = 8'h00; 
    ram[3896] = 8'h00; ram[3897] = 8'h00; ram[3898] = 8'h00; ram[3899] = 8'h00; 
    ram[3900] = 8'h00; ram[3901] = 8'h00; ram[3902] = 8'h00; ram[3903] = 8'h00; 
    ram[3904] = 8'h00; ram[3905] = 8'h00; ram[3906] = 8'h00; ram[3907] = 8'h00; 
    ram[3908] = 8'h00; ram[3909] = 8'h00; ram[3910] = 8'h00; ram[3911] = 8'h00; 
    ram[3912] = 8'h00; ram[3913] = 8'h00; ram[3914] = 8'h00; ram[3915] = 8'h00; 
    ram[3916] = 8'h00; ram[3917] = 8'h00; ram[3918] = 8'h00; ram[3919] = 8'h00; 
    ram[3920] = 8'h00; ram[3921] = 8'h00; ram[3922] = 8'h00; ram[3923] = 8'h00; 
    ram[3924] = 8'h00; ram[3925] = 8'h00; ram[3926] = 8'h00; ram[3927] = 8'h00; 
    ram[3928] = 8'h00; ram[3929] = 8'h00; ram[3930] = 8'h00; ram[3931] = 8'h00; 
    ram[3932] = 8'h00; ram[3933] = 8'h00; ram[3934] = 8'h00; ram[3935] = 8'h00; 
    ram[3936] = 8'h00; ram[3937] = 8'h00; ram[3938] = 8'h00; ram[3939] = 8'h00; 
    ram[3940] = 8'h00; ram[3941] = 8'h00; ram[3942] = 8'h00; ram[3943] = 8'h00; 
    ram[3944] = 8'h00; ram[3945] = 8'h00; ram[3946] = 8'h00; ram[3947] = 8'h00; 
    ram[3948] = 8'h00; ram[3949] = 8'h00; ram[3950] = 8'h00; ram[3951] = 8'h00; 
    ram[3952] = 8'h00; ram[3953] = 8'h00; ram[3954] = 8'h00; ram[3955] = 8'h00; 
    ram[3956] = 8'h00; ram[3957] = 8'h00; ram[3958] = 8'h00; ram[3959] = 8'h00; 
    ram[3960] = 8'h00; ram[3961] = 8'h00; ram[3962] = 8'h00; ram[3963] = 8'h00; 
    ram[3964] = 8'h00; ram[3965] = 8'h00; ram[3966] = 8'h00; ram[3967] = 8'h00; 
    ram[3968] = 8'h00; ram[3969] = 8'h00; ram[3970] = 8'h00; ram[3971] = 8'h00; 
    ram[3972] = 8'h00; ram[3973] = 8'h00; ram[3974] = 8'h00; ram[3975] = 8'h00; 
    ram[3976] = 8'h00; ram[3977] = 8'h00; ram[3978] = 8'h00; ram[3979] = 8'h00; 
    ram[3980] = 8'h00; ram[3981] = 8'h00; ram[3982] = 8'h00; ram[3983] = 8'h00; 
    ram[3984] = 8'h00; ram[3985] = 8'h00; ram[3986] = 8'h00; ram[3987] = 8'h00; 
    ram[3988] = 8'h00; ram[3989] = 8'h00; ram[3990] = 8'h00; ram[3991] = 8'h00; 
    ram[3992] = 8'h00; ram[3993] = 8'h00; ram[3994] = 8'h00; ram[3995] = 8'h00; 
    ram[3996] = 8'h00; ram[3997] = 8'h00; ram[3998] = 8'h00; ram[3999] = 8'h00; 
    ram[4000] = 8'h00; ram[4001] = 8'h00; ram[4002] = 8'h00; ram[4003] = 8'h00; 
    ram[4004] = 8'h00; ram[4005] = 8'h00; ram[4006] = 8'h00; ram[4007] = 8'h00; 
    ram[4008] = 8'h00; ram[4009] = 8'h00; ram[4010] = 8'h00; ram[4011] = 8'h00; 
    ram[4012] = 8'h00; ram[4013] = 8'h00; ram[4014] = 8'h00; ram[4015] = 8'h00; 
    ram[4016] = 8'h00; ram[4017] = 8'h00; ram[4018] = 8'h00; ram[4019] = 8'h00; 
    ram[4020] = 8'h00; ram[4021] = 8'h00; ram[4022] = 8'h00; ram[4023] = 8'h00; 
    ram[4024] = 8'h00; ram[4025] = 8'h00; ram[4026] = 8'h00; ram[4027] = 8'h00; 
    ram[4028] = 8'h00; ram[4029] = 8'h00; ram[4030] = 8'h00; ram[4031] = 8'h00; 
    ram[4032] = 8'h00; ram[4033] = 8'h00; ram[4034] = 8'h00; ram[4035] = 8'h00; 
    ram[4036] = 8'h00; ram[4037] = 8'h00; ram[4038] = 8'h00; ram[4039] = 8'h00; 
    ram[4040] = 8'h00; ram[4041] = 8'h00; ram[4042] = 8'h00; ram[4043] = 8'h00; 
    ram[4044] = 8'h00; ram[4045] = 8'h00; ram[4046] = 8'h00; ram[4047] = 8'h00; 
    ram[4048] = 8'h00; ram[4049] = 8'h00; ram[4050] = 8'h00; ram[4051] = 8'h00; 
    ram[4052] = 8'h00; ram[4053] = 8'h00; ram[4054] = 8'h00; ram[4055] = 8'h00; 
    ram[4056] = 8'h00; ram[4057] = 8'h00; ram[4058] = 8'h00; ram[4059] = 8'h00; 
    ram[4060] = 8'h00; ram[4061] = 8'h00; ram[4062] = 8'h00; ram[4063] = 8'h00; 
    ram[4064] = 8'h00; ram[4065] = 8'h00; ram[4066] = 8'h00; ram[4067] = 8'h00; 
    ram[4068] = 8'h00; ram[4069] = 8'h00; ram[4070] = 8'h00; ram[4071] = 8'h00; 
    ram[4072] = 8'h00; ram[4073] = 8'h00; ram[4074] = 8'h00; ram[4075] = 8'h00; 
    ram[4076] = 8'h00; ram[4077] = 8'h00; ram[4078] = 8'h00; ram[4079] = 8'h00; 
    ram[4080] = 8'h00; ram[4081] = 8'h00; ram[4082] = 8'h00; ram[4083] = 8'h00; 
    ram[4084] = 8'h00; ram[4085] = 8'h00; ram[4086] = 8'h00; ram[4087] = 8'h00; 
    ram[4088] = 8'h00; ram[4089] = 8'h00; ram[4090] = 8'h00; ram[4091] = 8'h00; 
    ram[4092] = 8'h00; ram[4093] = 8'h00; ram[4094] = 8'h00; ram[4095] = 8'h00; 
end

//-----------------------------------------------------------------------------
always @(posedge clk)
begin
    if (we)
        ram[addr] <= din;
    dout <= ram[addr];
end

endmodule
//-----------------------------------------------------------------------------
