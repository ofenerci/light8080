library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity c2sb_cpm_rom is
    port ( 
				clk						: in std_logic;
				addr					: in std_logic_vector(15 downto 0);
				data_out			: out std_logic_vector(7 downto 0)
		);
end c2sb_cpm_rom;

architecture internal of c2sb_cpm_rom is

signal rom_addr :         std_logic_vector(10 downto 0);
type t_rom is array(0 to 2047) of std_logic_vector(7 downto 0);

signal rom : t_rom := (

X"31",X"ff",X"3f",X"c3",X"40",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"c3",X"a5",X"07",X"00",X"00",X"00",X"00",X"00",
X"01",X"00",X"08",X"21",X"00",X"00",X"7e",X"77",
X"23",X"0b",X"78",X"b1",X"c2",X"46",X"00",X"cd",
X"f1",X"01",X"cd",X"18",X"02",X"21",X"f0",X"00",
X"cd",X"aa",X"02",X"cd",X"38",X"04",X"b7",X"c2",
X"d4",X"00",X"21",X"9a",X"06",X"cd",X"34",X"07",
X"21",X"1d",X"01",X"cd",X"aa",X"02",X"21",X"11",
X"43",X"cd",X"aa",X"02",X"21",X"36",X"01",X"cd",
X"aa",X"02",X"21",X"e1",X"00",X"11",X"1d",X"43",
X"06",X"0b",X"cd",X"99",X"02",X"21",X"89",X"06",
X"cd",X"34",X"07",X"3a",X"ef",X"42",X"b7",X"c2",
X"bb",X"00",X"cd",X"50",X"06",X"21",X"bf",X"01",
X"cd",X"aa",X"02",X"21",X"e1",X"00",X"cd",X"aa",
X"02",X"21",X"d4",X"01",X"cd",X"aa",X"02",X"cd",
X"19",X"02",X"cd",X"c2",X"02",X"21",X"df",X"01",
X"cd",X"aa",X"02",X"3e",X"01",X"d3",X"22",X"c3",
X"00",X"f2",X"76",X"21",X"a0",X"01",X"cd",X"aa",
X"02",X"21",X"e1",X"00",X"cd",X"aa",X"02",X"21",
X"ac",X"01",X"cd",X"aa",X"02",X"21",X"85",X"01",
X"cd",X"aa",X"02",X"76",X"21",X"3e",X"01",X"cd",
X"aa",X"02",X"21",X"85",X"01",X"cd",X"aa",X"02",
X"76",X"53",X"44",X"42",X"49",X"4f",X"53",X"20",
X"20",X"48",X"45",X"58",X"00",X"1b",X"63",X"00",
X"0a",X"1b",X"5b",X"33",X"36",X"6d",X"53",X"44",
X"2d",X"43",X"61",X"72",X"64",X"20",X"43",X"50",
X"2f",X"4d",X"20",X"62",X"6f",X"6f",X"74",X"6c",
X"6f",X"61",X"64",X"65",X"72",X"20",X"28",X"30",
X"2e",X"30",X"2e",X"31",X"29",X"0a",X"0d",X"0a",
X"1b",X"5b",X"30",X"6d",X"00",X"55",X"73",X"69",
X"6e",X"67",X"20",X"46",X"41",X"54",X"31",X"36",
X"20",X"76",X"6f",X"6c",X"75",X"6d",X"65",X"20",
X"1b",X"5b",X"33",X"35",X"6d",X"00",X"1b",X"5b",
X"30",X"6d",X"0a",X"0a",X"0d",X"00",X"0a",X"53",
X"44",X"20",X"63",X"61",X"72",X"64",X"20",X"6e",
X"6f",X"74",X"20",X"66",X"6f",X"75",X"6e",X"64",
X"20",X"6f",X"72",X"20",X"66",X"6f",X"72",X"6d",
X"61",X"74",X"20",X"69",X"73",X"20",X"6e",X"6f",
X"74",X"20",X"46",X"41",X"54",X"20",X"31",X"36",
X"3b",X"20",X"6e",X"6f",X"20",X"66",X"69",X"6c",
X"65",X"73",X"79",X"73",X"74",X"65",X"6d",X"20",
X"61",X"76",X"61",X"69",X"6c",X"61",X"62",X"6c",
X"65",X"2e",X"0a",X"0d",X"00",X"0a",X"1b",X"5b",
X"33",X"31",X"6d",X"53",X"79",X"73",X"74",X"65",
X"6d",X"20",X"68",X"61",X"6c",X"74",X"65",X"64",
X"2e",X"0a",X"0d",X"1b",X"5b",X"30",X"6d",X"00",
X"46",X"69",X"6c",X"65",X"20",X"27",X"1b",X"5b",
X"33",X"35",X"6d",X"00",X"1b",X"5b",X"30",X"6d",
X"27",X"20",X"6e",X"6f",X"74",X"20",X"66",X"6f",
X"75",X"6e",X"64",X"2e",X"0a",X"0d",X"00",X"0a",
X"4c",X"6f",X"61",X"64",X"69",X"6e",X"67",X"20",
X"66",X"69",X"6c",X"65",X"20",X"27",X"1b",X"5b",
X"33",X"35",X"6d",X"00",X"1b",X"5b",X"30",X"6d",
X"27",X"2e",X"2e",X"2e",X"20",X"20",X"00",X"68",
X"20",X"62",X"79",X"74",X"65",X"73",X"20",X"6c",
X"6f",X"61",X"64",X"65",X"64",X"2e",X"0a",X"0d",
X"00",X"c9",X"21",X"ff",X"01",X"cd",X"aa",X"02",
X"21",X"85",X"01",X"cd",X"aa",X"02",X"76",X"1b",
X"5b",X"33",X"33",X"6d",X"50",X"4f",X"53",X"54",
X"20",X"66",X"61",X"69",X"6c",X"75",X"72",X"65",
X"2e",X"0a",X"0d",X"1b",X"5b",X"30",X"6d",X"00",
X"c9",X"21",X"00",X"00",X"e5",X"cd",X"b1",X"03",
X"b7",X"ca",X"2f",X"02",X"cd",X"31",X"02",X"e1",
X"4f",X"af",X"47",X"09",X"c3",X"1c",X"02",X"e1",
X"c9",X"21",X"00",X"40",X"7e",X"23",X"fe",X"3a",
X"c2",X"77",X"02",X"cd",X"18",X"03",X"32",X"c6",
X"40",X"cd",X"18",X"03",X"32",X"c8",X"40",X"cd",
X"18",X"03",X"32",X"c7",X"40",X"cd",X"18",X"03",
X"fe",X"00",X"c2",X"72",X"02",X"3a",X"c7",X"40",
X"5f",X"3a",X"c8",X"40",X"57",X"3a",X"c6",X"40",
X"4f",X"c5",X"d5",X"cd",X"18",X"03",X"d1",X"c1",
X"12",X"13",X"0d",X"c2",X"61",X"02",X"3a",X"c6",
X"40",X"c9",X"fe",X"01",X"c2",X"77",X"02",X"af",
X"c9",X"1a",X"b7",X"c8",X"be",X"c0",X"23",X"13",
X"0d",X"c8",X"c3",X"79",X"02",X"7e",X"12",X"23",
X"13",X"0b",X"78",X"b1",X"c2",X"85",X"02",X"c9",
X"12",X"13",X"0b",X"78",X"b1",X"c2",X"90",X"02",
X"c9",X"05",X"7e",X"fe",X"00",X"ca",X"a7",X"02",
X"23",X"12",X"13",X"05",X"c2",X"9a",X"02",X"af",
X"12",X"c9",X"4e",X"79",X"b7",X"c8",X"23",X"e5",
X"cd",X"2a",X"04",X"e1",X"c3",X"aa",X"02",X"0e",
X"0d",X"cd",X"2a",X"04",X"0e",X"0a",X"cd",X"2a",
X"04",X"c9",X"7c",X"e5",X"cd",X"cd",X"02",X"e1",
X"7d",X"cd",X"cd",X"02",X"c9",X"f5",X"0f",X"0f",
X"0f",X"0f",X"cd",X"da",X"02",X"f1",X"cd",X"da",
X"02",X"c9",X"e6",X"0f",X"21",X"e8",X"02",X"4f",
X"06",X"00",X"09",X"4e",X"cd",X"2a",X"04",X"c9",
X"30",X"31",X"32",X"33",X"34",X"35",X"36",X"37",
X"38",X"39",X"61",X"62",X"63",X"64",X"65",X"66",
X"f6",X"20",X"fe",X"30",X"da",X"16",X"03",X"fe",
X"3a",X"d2",X"07",X"03",X"d6",X"30",X"c9",X"fe",
X"61",X"da",X"16",X"03",X"fe",X"67",X"d2",X"16",
X"03",X"d6",X"61",X"c6",X"0a",X"c9",X"37",X"c9",
X"7e",X"23",X"e5",X"cd",X"f8",X"02",X"e1",X"07",
X"07",X"07",X"07",X"e6",X"f0",X"47",X"7e",X"23",
X"e5",X"cd",X"f8",X"02",X"e1",X"e6",X"0f",X"b0",
X"c9",X"22",X"c4",X"40",X"c5",X"e5",X"7c",X"cd",
X"cd",X"02",X"e1",X"e5",X"7d",X"cd",X"cd",X"02",
X"0e",X"3a",X"cd",X"2a",X"04",X"0e",X"20",X"cd",
X"2a",X"04",X"e1",X"c1",X"0e",X"10",X"7e",X"e5",
X"c5",X"cd",X"cd",X"02",X"0e",X"20",X"cd",X"2a",
X"04",X"c1",X"c5",X"79",X"fe",X"09",X"c2",X"66",
X"03",X"0e",X"20",X"cd",X"2a",X"04",X"c1",X"e1",
X"23",X"0d",X"c2",X"4e",X"03",X"0e",X"10",X"e5",
X"c5",X"0e",X"7c",X"cd",X"2a",X"04",X"0e",X"20",
X"cd",X"2a",X"04",X"0e",X"20",X"cd",X"2a",X"04",
X"2a",X"c4",X"40",X"06",X"10",X"7e",X"23",X"e5",
X"c5",X"57",X"e6",X"80",X"c2",X"95",X"03",X"7a",
X"e6",X"f0",X"c2",X"9d",X"03",X"0e",X"2e",X"cd",
X"2a",X"04",X"c3",X"a1",X"03",X"4a",X"cd",X"2a",
X"04",X"c1",X"e1",X"05",X"c2",X"85",X"03",X"cd",
X"b7",X"02",X"c1",X"e1",X"05",X"c2",X"31",X"03",
X"c9",X"0e",X"00",X"21",X"00",X"40",X"e5",X"c5",
X"cd",X"d0",X"03",X"c1",X"e1",X"b7",X"ca",X"cc",
X"03",X"0c",X"77",X"23",X"fe",X"0a",X"ca",X"cc",
X"03",X"c3",X"b6",X"03",X"af",X"77",X"79",X"c9",
X"2a",X"35",X"43",X"7c",X"e6",X"fe",X"c2",X"0c",
X"04",X"3a",X"39",X"43",X"bd",X"c2",X"f8",X"03",
X"3a",X"3a",X"43",X"bc",X"c2",X"f8",X"03",X"2a",
X"33",X"43",X"3a",X"37",X"43",X"bd",X"c2",X"f8",
X"03",X"3a",X"37",X"43",X"bc",X"ca",X"12",X"04",
X"af",X"32",X"ef",X"42",X"2a",X"35",X"43",X"01",
X"d9",X"40",X"09",X"7e",X"2a",X"35",X"43",X"23",
X"22",X"35",X"43",X"c9",X"cd",X"78",X"06",X"c3",
X"f8",X"03",X"3e",X"02",X"32",X"ef",X"42",X"af",
X"c9",X"db",X"20",X"e6",X"01",X"ca",X"22",X"04",
X"af",X"c9",X"3e",X"ff",X"c9",X"db",X"21",X"e6",
X"7f",X"c9",X"db",X"20",X"2f",X"e6",X"80",X"ca",
X"2a",X"04",X"79",X"e6",X"7f",X"d3",X"21",X"c9",
X"d3",X"93",X"d3",X"95",X"06",X"14",X"3e",X"ff",
X"32",X"c9",X"40",X"c5",X"cd",X"06",X"05",X"c1",
X"05",X"c2",X"3e",X"04",X"d3",X"94",X"0e",X"00",
X"cd",X"44",X"05",X"3a",X"d1",X"40",X"e6",X"80",
X"c2",X"03",X"05",X"0e",X"01",X"cd",X"44",X"05",
X"3a",X"d1",X"40",X"e6",X"01",X"c2",X"5b",X"04",
X"21",X"00",X"00",X"22",X"eb",X"42",X"22",X"ed",
X"42",X"cd",X"7a",X"07",X"2a",X"d7",X"42",X"7c",
X"fe",X"aa",X"c2",X"fd",X"04",X"7d",X"fe",X"55",
X"c2",X"fd",X"04",X"3a",X"9b",X"42",X"fe",X"06",
X"c2",X"00",X"05",X"2a",X"9f",X"42",X"22",X"e7",
X"42",X"2a",X"e7",X"42",X"22",X"eb",X"42",X"21",
X"00",X"00",X"22",X"ed",X"42",X"cd",X"7a",X"07",
X"21",X"04",X"41",X"11",X"11",X"43",X"06",X"0c",
X"cd",X"99",X"02",X"2a",X"ea",X"40",X"22",X"e9",
X"42",X"3a",X"e6",X"40",X"32",X"10",X"43",X"2a",
X"e7",X"40",X"44",X"4d",X"2a",X"e7",X"42",X"09",
X"22",X"2b",X"43",X"e5",X"2a",X"ef",X"40",X"22",
X"29",X"43",X"44",X"4d",X"09",X"44",X"4d",X"e1",
X"09",X"22",X"2d",X"43",X"2a",X"e9",X"42",X"7d",
X"0f",X"0f",X"0f",X"0f",X"e6",X"0f",X"4f",X"7c",
X"07",X"07",X"07",X"07",X"e6",X"f0",X"b1",X"4f",
X"7c",X"0f",X"0f",X"0f",X"0f",X"e6",X"0f",X"47",
X"4d",X"01",X"20",X"00",X"2a",X"2d",X"43",X"09",
X"22",X"2f",X"43",X"af",X"c9",X"3e",X"01",X"c9",
X"3e",X"02",X"c9",X"3e",X"04",X"c9",X"1e",X"08",
X"3a",X"c9",X"40",X"17",X"32",X"c9",X"40",X"da",
X"17",X"05",X"d3",X"90",X"c3",X"19",X"05",X"d3",
X"91",X"d3",X"92",X"00",X"d3",X"93",X"db",X"88",
X"17",X"3a",X"ca",X"40",X"17",X"32",X"ca",X"40",
X"00",X"1d",X"c2",X"08",X"05",X"3a",X"ca",X"40",
X"c9",X"7e",X"23",X"e5",X"c5",X"32",X"c9",X"40",
X"cd",X"06",X"05",X"c1",X"e1",X"0b",X"78",X"b1",
X"c2",X"31",X"05",X"c9",X"21",X"cb",X"40",X"79",
X"77",X"23",X"af",X"06",X"05",X"77",X"23",X"05",
X"c2",X"4d",X"05",X"79",X"fe",X"00",X"c2",X"61",
X"05",X"3e",X"94",X"32",X"d0",X"40",X"c3",X"9d",
X"05",X"fe",X"10",X"c2",X"6e",X"05",X"3e",X"02",
X"32",X"ce",X"40",X"c3",X"9d",X"05",X"fe",X"51",
X"c2",X"8d",X"05",X"21",X"eb",X"42",X"37",X"3f",
X"7e",X"23",X"17",X"32",X"ce",X"40",X"7e",X"23",
X"17",X"32",X"cd",X"40",X"7e",X"23",X"17",X"32",
X"cc",X"40",X"c3",X"9d",X"05",X"fe",X"01",X"c2",
X"95",X"05",X"c3",X"9d",X"05",X"fe",X"3a",X"c2",
X"9d",X"05",X"c3",X"9d",X"05",X"21",X"cb",X"40",
X"7e",X"e6",X"3f",X"f6",X"40",X"77",X"21",X"d0",
X"40",X"7e",X"f6",X"01",X"77",X"21",X"cb",X"40",
X"01",X"06",X"00",X"cd",X"31",X"05",X"cd",X"c5",
X"05",X"32",X"d1",X"40",X"b7",X"c2",X"c2",X"05",
X"af",X"c9",X"af",X"3c",X"c9",X"21",X"64",X"00",
X"22",X"d7",X"40",X"3e",X"ff",X"32",X"c9",X"40",
X"cd",X"06",X"05",X"3a",X"ca",X"40",X"fe",X"ff",
X"c0",X"2a",X"d7",X"40",X"2b",X"22",X"d7",X"40",
X"7c",X"b5",X"c2",X"cb",X"05",X"3e",X"ff",X"c9",
X"11",X"3f",X"43",X"21",X"43",X"43",X"37",X"3f",
X"cd",X"fd",X"05",X"cd",X"fd",X"05",X"cd",X"fd",
X"05",X"cd",X"fd",X"05",X"c9",X"1a",X"8e",X"12",
X"23",X"13",X"c9",X"21",X"00",X"00",X"22",X"41",
X"43",X"22",X"3f",X"43",X"22",X"45",X"43",X"2a",
X"31",X"43",X"2b",X"2b",X"22",X"43",X"43",X"3a",
X"10",X"43",X"47",X"cd",X"e8",X"05",X"05",X"c2",
X"1b",X"06",X"2a",X"2f",X"43",X"22",X"43",X"43",
X"21",X"00",X"00",X"22",X"45",X"43",X"cd",X"e8",
X"05",X"2a",X"33",X"43",X"22",X"43",X"43",X"21",
X"00",X"00",X"22",X"45",X"43",X"cd",X"e8",X"05",
X"2a",X"3f",X"43",X"22",X"eb",X"42",X"2a",X"41",
X"43",X"22",X"ed",X"42",X"cd",X"7a",X"07",X"c9",
X"2a",X"0a",X"43",X"22",X"31",X"43",X"af",X"6f",
X"67",X"22",X"35",X"43",X"22",X"33",X"43",X"2a",
X"0c",X"43",X"44",X"7c",X"e6",X"01",X"67",X"22",
X"39",X"43",X"78",X"0f",X"e6",X"7f",X"6f",X"26",
X"00",X"22",X"37",X"43",X"cd",X"03",X"06",X"c9",
X"2a",X"33",X"43",X"23",X"22",X"33",X"43",X"21",
X"00",X"00",X"22",X"35",X"43",X"cd",X"03",X"06",
X"c9",X"11",X"1d",X"43",X"21",X"f0",X"42",X"0e",
X"0b",X"cd",X"79",X"02",X"c0",X"af",X"32",X"ef",
X"42",X"c9",X"3a",X"fb",X"42",X"6f",X"fe",X"0f",
X"ca",X"a8",X"06",X"e6",X"08",X"c2",X"ab",X"06",
X"af",X"3c",X"c9",X"21",X"f0",X"42",X"11",X"11",
X"43",X"06",X"0c",X"cd",X"99",X"02",X"af",X"c9",
X"3a",X"fb",X"42",X"6f",X"fe",X"0f",X"c8",X"e6",
X"08",X"c2",X"f0",X"06",X"7d",X"e6",X"10",X"c2",
X"d3",X"06",X"21",X"f3",X"06",X"cd",X"aa",X"02",
X"c3",X"d9",X"06",X"21",X"f9",X"06",X"cd",X"aa",
X"02",X"21",X"f0",X"42",X"06",X"0c",X"11",X"80",
X"40",X"cd",X"99",X"02",X"21",X"80",X"40",X"cd",
X"aa",X"02",X"21",X"ff",X"06",X"cd",X"aa",X"02",
X"af",X"3c",X"c9",X"1b",X"5b",X"33",X"35",X"6d",
X"00",X"1b",X"5b",X"33",X"34",X"6d",X"00",X"1b",
X"5b",X"30",X"6d",X"0a",X"0d",X"00",X"21",X"d9",
X"40",X"0e",X"10",X"7e",X"fe",X"e5",X"ca",X"25",
X"07",X"fe",X"00",X"c8",X"e5",X"c5",X"11",X"f0",
X"42",X"01",X"20",X"00",X"cd",X"85",X"02",X"cd",
X"30",X"07",X"c1",X"e1",X"c8",X"11",X"20",X"00",
X"19",X"0d",X"c2",X"0b",X"07",X"af",X"3c",X"c9",
X"2a",X"e5",X"42",X"e9",X"22",X"e5",X"42",X"3e",
X"01",X"32",X"ef",X"42",X"2a",X"2d",X"43",X"22",
X"eb",X"42",X"21",X"00",X"00",X"22",X"ed",X"42",
X"cd",X"7a",X"07",X"2a",X"e9",X"42",X"e5",X"cd",
X"06",X"07",X"e1",X"c8",X"7d",X"d6",X"10",X"6f",
X"7c",X"de",X"00",X"b5",X"c8",X"e5",X"cd",X"64",
X"07",X"c3",X"4f",X"07",X"2a",X"eb",X"42",X"23",
X"22",X"eb",X"42",X"7c",X"b5",X"c2",X"7a",X"07",
X"2a",X"ed",X"42",X"23",X"22",X"ed",X"42",X"c3",
X"7a",X"07",X"0e",X"51",X"cd",X"44",X"05",X"cd",
X"c5",X"05",X"fe",X"fe",X"c2",X"7f",X"07",X"21",
X"d9",X"40",X"01",X"02",X"02",X"e5",X"c5",X"3e",
X"ff",X"32",X"c9",X"40",X"cd",X"06",X"05",X"3a",
X"ca",X"40",X"c1",X"e1",X"77",X"23",X"0b",X"78",
X"b1",X"c2",X"8d",X"07",X"c9",X"22",X"3d",X"43",
X"e1",X"e5",X"22",X"3b",X"43",X"2a",X"3d",X"43",
X"f5",X"d5",X"e5",X"c5",X"21",X"cc",X"07",X"cd",
X"aa",X"02",X"2a",X"3b",X"43",X"cd",X"c2",X"02",
X"21",X"d0",X"07",X"cd",X"aa",X"02",X"c1",X"e1",
X"d1",X"f1",X"fb",X"c9",X"50",X"43",X"3d",X"00",
X"0a",X"0d",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"

);


begin


-- Program memory (it's RAM really)
rom_addr <= addr(10 downto 0);
process(clk)
begin
  if (clk'event and clk='1') then
    data_out <= rom(conv_integer(rom_addr));
  end if;
end process;

end internal;
